module pspoltop ( SCLK, CRST, WRST, ADS, WR, RDYOL, RDYOLCNT, IBSY, PA02, PA, 
    BE, CA, PDH, PDLIN, PDLOUT, PDCNT, CDIN, CDOUT, CDCNT, LIN, LOUT, LCNT, 
    CPIN, CPOUT, LPIN, LPOUT, CRCE, CRWE, CROE, LRQ, LGR, LASIN, LASOUT, LWR, 
    LDS, LDK, LDL0, LPDIN, LPDOUT, LTC0, LCMDCNT, LPDCNT, LBSY, LBER, SWIT, 
    DTFL, HINT, phtri );
input  [31:3] PA;
output [3:0] CPOUT;
input  [7:0] BE;
input  [31:0] PDLIN;
input  [59:0] CDIN;
input  [31:0] LIN;
output [18:0] CA;
output [63:32] PDH;
output [31:0] LOUT;
input  [3:0] CPIN;
output [31:0] PDLOUT;
output [59:0] CDOUT;
input  [3:0] LPIN;
output [3:0] LPOUT;
input  SCLK, CRST, WRST, ADS, WR, IBSY, PA02, LGR, LASIN, LDK, LPDIN, LBSY, 
    LBER, SWIT, DTFL, HINT, phtri;
output RDYOL, RDYOLCNT, PDCNT, CDCNT, LCNT, CRCE, CRWE, CROE, LRQ, LASOUT, LWR, 
    LDS, LDL0, LPDOUT, LTC0, LCMDCNT, LPDCNT;
    wire \SADR/operand[7] , \SADR/operand[26] , \stream3[7] , \pk_dpr_h[14] , 
        \pk_sra1_h[8] , \pk_idcw_h[1] , \REGF/RI_DPR[1] , \ADOSEL/n4132 , 
        \CODEIF/n4031 , \CODEQ/nqueue1[31] , \CODEQ/nqueue1[28] , eaccbsel, 
        \LBUS/n1393 , \LBUS/n1412 , ph_srcadr2_h, \SADR/pgaddwx[6] , 
        \pk_scdl_h[25] , \pk_scdl_h[16] , \REGF/n8244 , pkaluopc, 
        \pgbluext[5] , \CONS/SACO[10] , \BLU/n1478 , \PDOSEL/n107 , 
        \REGF/n8174 , \SADR/pgaddwyz[1] , \pk_indz_h[18] , \pk_s1ba_h[0] , 
        \pk_scdl_h[6] , \REGF/n8153 , \pkdptout[15] , \pk_sefl_h[14] , 
        \pgmuxout[27] , \pgaluina[17] , \CODEQ/nqueue2[58] , 
        \CODEQ/nqueue2[41] , \SADR/sadr[18] , \pk_s6ba_h[14] , \pk_s01l_h[3] , 
        ph_pccons_h, \ADOSEL/n4115 , \CODEIF/n4016 , \pk_s45l_h[18] , 
        \pk_sefl_h[27] , \REGF/RO_ACC[8] , \pgmuxout[14] , \pgaluina[24] , 
        \LBUS/n1435 , cif_byte, \LDIS/ldexcl[2] , \pkdptout[26] , 
        \CODEIF/n3866 , \PDOSEL/n120 , \pk_stdat[13] , \LDIS/n3129 , 
        \CONS/n601 , \BLU/n1563 , \REGF/RO_EACC[0] , \pgaluinb[9] , 
        \CONS/n531 , \MAIN/n3624 , \pk_s23l_h[4] , \pk_stdat[20] , 
        \pk_scba_h[1] , \pk_rread_h[10] , \pk_s67l_h[24] , \pk_s67l_h[17] , 
        \REGF/RO_PCON[22] , \pk_rwrit_h[43] , \pk_rread_h[23] , \stream2[25] , 
        \BLU/n1544 , \CONS/n626 , \pk_pcs1_h[8] , \SADR/pgaddwxy[8] , 
        \pk_scba_h[13] , \REGF/RI_PCOH[3] , \REGF/RO_PCON[11] , 
        \pk_idcx_h[14] , wdpr, \CONS/n578 , \pgsdprlh[3] , \pk_saseo_h[0] , 
        \LDCHK/n3249 , \pk_s23l_h[22] , \pk_s23l_h[11] , \CODEIF/n3883 , 
        \CODEIF/n3913 , \LDIS/n3160 , \CONS/n648 , \REG_2/ncnt2[1] , 
        \pk_idcy_h[3] , \REG_2/ncnt1[2] , \LDIS/n3147 , \SADR/operand[15] , 
        \pk_s45l_h[6] , \CODEIF/n3934 , \CODEIF/pfctr415[17] , \ALUIS/n3679 , 
        \pk_indz_h[5] , \REGF/n8191 , \pk_s0ba_h[7] , ph_ldaoutenh3, 
        \SAEXE/*cell*3651/U4/CONTROL1 , n10734, \stream3[26] , \stream3[15] , 
        \pk_spr_h[7] , \SADR/pgaddxz[21] , \SADR/pgaddwxy[14] , 
        \pgregadrh[11] , \pk_s89l_h[0] , ph_sacons_h, \pk_adb_h[6] , ph_selldl, 
        \pk_s67l_h[1] , \pk_sabl_h[21] , \pk_idcy_h[19] , \ALUIS/n3745 , 
        \pk_sabl_h[12] , \REGF/RI_SPR[4] , \pgregadrh[22] , 
        \CODEIF/pfctr415[2] , \CODEIF/n3998 , \pgsdprlh[11] , 
        \REGF/RO_LLPSAS[15] , \CODEIF/fddacnt_in , \PDOSEL/n98 , 
        \SADR/pgaddxz[12] , \pk_s89l_h[18] , \pk_saco_lh[0] , ph_lbend, 
        \BLU/n1586 , \stream4[44] , \pgsdprlh[22] , \pk_s5ba_h[15] , 
        \pk_sbba_h[6] , \REGF/RO_ERFA[0] , \REGF/n8091 , \REGF/n8101 , 
        \pk_sra2_h[15] , \pk_s5ba_h[2] , \LBUS/*cell*3982/U119/CONTROL1 , 
        \REGF/n8231 , \pk_trba_h[7] , \SADR/pgaddwxy[1] , \SADR/pgaddwxz[2] , 
        \pk_s1ba_h[11] , \pk_s8ba_h[17] , \CODEIF/n4044 , \pk_rread_h[5] , 
        \ADOSEL/n4147 , \pk_s23l_h[18] , \LBUS/n1440 , \CONS/n748 , 
        \REGF/RI_SRA12M[25] , \REGF/n8216 , \CODEIF/n3983 , 
        \MAIN/excep_enable , \PDOSEL/n155 , \REGF/RO_ACC[15] , 
        \ALUSHT/pkshtout[7] , phrelbwrh, \pgsadrh[7] , \REGF/RI_SRA12M[16] , 
        \REGF/n8126 , \REGF/RO_PSTA[17] , \pgfdout[1] , \ALUSHT/pkaluout[2] , 
        \REGF/RO_ACC[26] , \CODEIF/pgctrinc[13] , \REGF/RO_LPSAS2156[2] , 
        \pgsadrh[21] , \pgsadrh[12] , \pk_s89l_h[22] , \pk_stdat[2] , 
        \REGF/pk_idcy_h[27] , \SAEXE/n434 , \pkbludgh[7] , \LDCHK/n3275 , 
        \MAIN/WP_PC , \MAIN/*cell*4603/U16/CONTROL1 , \pgld32[14] , 
        \LBUS/*cell*3982/U148/CONTROL1 , \CONS/n544 , \pgsdprlh[18] , 
        \pk_idcw_h[14] , po_imdselh, \ALUIS/n3662 , \BLU/n1516 , 
        \SADR/operand[3] , \SADR/pgaddwz[16] , \pgregadrh[18] , 
        \SADR/segbase[13] , \pk_s89l_h[11] , \pk_saco_lh[9] , \BLU/n1486 , 
        \stream4[54] , \pgld32[27] , \CONS/n674 , \pk_s01l_h[24] , 
        \pk_s67l_h[8] , \pk_idcy_h[10] , \ALUIS/n3645 , \REGF/RI_SRDA[5] , 
        \pk_pcs1_h[15] , \CODEIF/n3898 , \CODEIF/n3908 , \pk_s01l_h[17] , 
        \pk_s89l_h[9] , \pk_sefl_h[3] , \pk_idcy_h[23] , \CONS/n653 , 
        \BLU/n1531 , \LDCHK/n3252 , \REGF/pk_s5ba_h[18] , \SAEXE/n413 , 
        \CONS/n563 , \pk_sabl_h[31] , \pk_sabl_h[28] , \pk_indz_h[22] , 
        \pk_sdba_h[16] , \REGF/pk_exco_h[0] , \pk_s45l_h[11] , \pk_psae_h[0] , 
        \pk_idcx_h[5] , \LDIS/n3115 , \SADR/sadr[11] , \pk_s4ba_h[5] , 
        \REGF/RO_ACC[1] , \CODEIF/n3966 , \pk_spr_h[3] , \pk_sra1_h[1] , 
        \pk_indz_h[11] , \SADR/sadr[22] , \pk_s1ba_h[9] , \REGF/pk_scti_h[6] , 
        \REGF/n8053 , \MAIN/n3618 , \pk_s45l_h[22] , \SADR/m_fadrl[8] , 
        \REGF/n8074 , \LBUS/n1605 , \CODEQ/nqueue2[51] , \CODEQ/nqueue1[12] , 
        \CODEQ/nqueue2[48] , \pk_idcw_h[8] , \REGF/RI_DPR[8] , 
        \CODEQ/nqueue1[38] , \CODEQ/nqueue1[21] , \SAEXE/relbwrh , 
        \SADR/pgaddyz[14] , \SADR/pgaddxyz[5] , \pk_sfba_h[4] , 
        \pk_rwrit_h[53] , \REGF/RO_ERRA[16] , \REGF/pk_indz_h[26] , 
        \CODEIF/n3941 , \LDIS/n3132 , \BLU/n1578 , \SAEXE/srcwrit , 
        \CONS/SACO[19] , \pk_pcs1_h[1] , \pk_rread_h[33] , ph_ixco_h, 
        \CONS/n726 , \MAIN/sw_end , \ALUIS/n3730 , \REGF/RO_PCON[18] , 
        \pk_rread_h[19] , \pk_scba_h[8] , \REGF/RO_ERRA[25] , \CONS/n586 , 
        \pk_rwrit_h[60] , \REGF/n8148 , \REGF/D2_HINT , \pgaluinb[0] , 
        \SADR/pgaddwyz[8] , \pk_adb_h[27] , \LBUS/*cell*3982/U71/CONTROL1 , 
        \pgaluina[3] , \LDCHK/n3290 , \SAEXE/trsc1_h , \SADR/pgovfwxy , 
        \pk_adb_h[14] , \LDCHK/n3300 , \pk_s2ba_h[10] , \LBUS/n1409 , 
        \LBUS/n1599 , \CONS/n691 , \CONS/n701 , \pk_sbba_h[2] , \pk_sabl_h[6] , 
        \REGF/RO_EACC[9] , \ALUIS/n3717 , \ADOSEL/n4129 , \ALUIS/n3687 , 
        pgiaendp, \pgsdprlh[15] , \pk_idcw_h[19] , \pk_saco_lh[4] , 
        \stream4[59] , \stream4[40] , \CONS/n734 , \PDOSEL/n129 , 
        \ALUIS/n3722 , \pgld32[19] , \CONS/n594 , \CMPX/n1051 , 
        \SADR/pgaddxz[16] , \pk_s5ba_h[11] , \SADR/pgaddwxy[23] , 
        \pgregadrh[15] , \pk_sabl_h[25] , \SADR/pgaddwxy[10] , \pk_s89l_h[4] , 
        \pk_adb_h[2] , \LDCHK/n3282 , \LDCHK/n3312 , \CODEIF/n3848 , 
        \CODEIF/pfctr415[6] , ph_pdhen_h, \CONS/n683 , \CONS/n713 , 
        \pk_s01l_h[30] , \pk_s01l_h[29] , \pk_sabl_h[16] , \REGF/RI_SPR[0] , 
        \BLU/n1471 , \pk_s67l_h[5] , \pk_pcs1_h[18] , \REGF/RI_SRDA[8] , 
        \SADR/operand[22] , \pk_sra2_h[18] , \SADR/lmtaddr[13] , 
        \CODEIF/n4038 , \ALUIS/n3695 , \pk_rread_h[8] , \ALUIS/n3705 , 
        \stream3[32] , \CODEIF/pfctr415[13] , \CODEIF/n3974 , 
        \SADR/operand[11] , \stream3[18] , \pk_s0ba_h[3] , 
        \REGF/pk_idcx_h[27] , \PDOSEL/n74 , \pk_indz_h[1] , \stream3[3] , 
        \pk_dpr_h[10] , \pk_scba_h[17] , \pk_s23l_h[26] , \pk_s45l_h[2] , 
        \REGF/pk_s1ba_h[18] , stage_b, \pgsdprlh[7] , \pk_scba_h[5] , 
        \pk_s23l_h[15] , \pk_idcx_h[10] , \pk_idcy_h[7] , \REGF/n8066 , 
        \CONS/n538 , po_opcsel_h, \REGF/RO_ACC[18] , \pk_s67l_h[13] , 
        \pk_idcx_h[23] , \CODEIF/n3953 , \LDIS/n3120 , \CONS/n608 , 
        \LDCHK/n3267 , \REGF/RO_PCON[26] , ph_dec_dh, \SAEXE/n426 , 
        \pk_rread_h[14] , \REGF/n8198 , \stream2[12] , \CONS/n556 , 
        \SADR/pgaddxyz[8] , \pk_sfba_h[9] , \REGF/RI_PCOH[7] , \CONS/n347 , 
        \REGF/RO_PCON[15] , \pk_dpr_h[23] , \pk_s67l_h[20] , \ALUIS/n3670 , 
        \pk_dpr_h[19] , \SADR/pgaddwx[2] , \SADR/pgaddyz[19] , 
        \SADR/pgaddwyz[5] , \pk_rwrit_h[47] , \pk_rread_h[27] , \stream2[21] , 
        \CONS/n666 , \BLU/n1494 , \pk_stdat[17] , \REGF/RO_EACC[4] , 
        \BLU/n1504 , \ALUIS/n3657 , \pk_adb_h[19] , \CONS/n641 , \BLU/n1523 , 
        \SAEXE/singlen , \pk_s23l_h[0] , \LDCHK/n3240 , \SAEXE/rf_srcadr2_h , 
        \SADR/m_fadrl[5] , \pk_s1ba_h[4] , \pk_sefl_h[10] , ph_ciwt_h, 
        write_pr_h, \CONS/n571 , \pgbluext[27] , \pgaluina[13] , 
        \CODEQ/nqueue2[45] , \pk_s4ba_h[8] , \pk_scdl_h[2] , \REGF/n8083 , 
        \REGF/n8113 , \pgmuxout[23] , \pkdptout[11] , \pkdptout[22] , 
        \REGF/n8223 , \pk_s6ba_h[10] , \pk_s01l_h[7] , \pk_sefl_h[23] , 
        \pk_idcx_h[8] , \pgmuxout[10] , \PDOSEL/n160 , \LDIS/ldexcl[6] , 
        \pgaluina[20] , \pk_scdl_h[12] , ph_baccwt_h, \ADOSEL/n4155 , 
        ph_bitsrc_h, \pk_idcw_h[5] , \REGF/n8204 , \pgbluext[1] , 
        \PDOSEL/n147 , \CODEIF/n3991 , \CONS/SACO[14] , \LBUS/n1452 , 
        \REGF/RI_DPR[5] , \CODEQ/nqueue1[35] , \SADR/pgaddyz[23] , 
        \SADR/pgaddyz[10] , \SADR/seglmterr , \pk_scdl_h[21] , \REGF/n8134 , 
        \pk_s23l_h[9] , \pk_adb_h[23] , po_ptrsel_h, \pgaluina[7] , 
        \pk_s2ba_h[14] , \pk_sabl_h[2] , ph_lbwrh, \pgaluinb[4] , \LBUS/n1449 , 
        \CONS/n741 , \REG_2/n410 , \pk_sfba_h[0] , \pk_adb_h[10] , 
        \pk_s67l_h[30] , \pk_s67l_h[29] , \pk_pcs1_h[5] , ph_srcsl_h, 
        \REGF/RO_ERRA[21] , \REGF/RO_ERRA[12] , \pk_rwrit_h[57] , 
        \pk_rread_h[37] , \REGF/n8238 , \pk_rwrit_h[64] , \REGF/n8108 , 
        \REGF/n8098 , \pk_sra1_h[5] , \SADR/pgaddxyz[1] , \pk_scdl_h[31] , 
        \pk_scdl_h[28] , \REGF/RO_TRCO[27] , \pgbluext[8] , 
        \CODEQ/nqueue1[16] , \CODEIF/n3891 , \CODEIF/n3901 , \BLU/n1538 , 
        \pk_indz_h[15] , \SADR/sadr[15] , \REGF/RO_ACC[5] , \pgmuxout[19] , 
        ph_exe_ch, \LBUS/n_2439 , \CODEQ/nqueue1[25] , \pk_s4ba_h[1] , 
        \CODEIF/n3926 , \pk_sdba_h[12] , \pk_s45l_h[15] , \LDIS/n3155 , 
        \pk_psae_h[4] , \pk_idcx_h[1] , \pgaluina[29] , \pgaluina[30] , 
        \pk_sefl_h[19] , \CODEQ/nqueue2[55] , \SADR/sadr[26] , \pk_s45l_h[26] , 
        \REGF/n8183 , \pkdptout[18] , \REGF/pk_scti_h[2] , \SADR/pgaddwz[21] , 
        \pk_s01l_h[20] , \REGF/RI_SPR[9] , \CONS/n613 , \BLU/n1571 , 
        \SADR/pgaddwz[12] , \SADR/pgaddwxy[19] , \SADR/segbase[17] , 
        \REGF/RI_SRDA[1] , \pk_pcs1_h[11] , \CODEIF/n3948 , \pk_idcy_h[14] , 
        \pk_s01l_h[13] , \pk_sefl_h[7] , \CONS/n523 , \SAEXE/srcwt_st , 
        \REGF/pk_idcw_h[27] , \SADR/operand[18] , \stream3[11] , 
        \pk_sra2_h[22] , \SADR/pgaddwxy[5] , \pgsadrh[25] , \pgsadrh[16] , 
        \pk_s89l_h[26] , \pk_stdat[6] , \pkbludgh[3] , \MAIN/n3611 , 
        \LDCHK/n3235 , \pgld32[10] , \pk_idcw_h[23] , \REGF/RO_LPSAS2156[6] , 
        \stream4[50] , \pgld32[23] , \CONS/n634 , \stream4[49] , \BLU/n1556 , 
        \pk_s8ba_h[13] , \pk_s89l_h[15] , \REGF/RI_SRA12M[21] , 
        \pk_idcw_h[10] , \MAIN/cstregw_inhibith , pk_pcser_h, \CODEIF/n4023 , 
        \REGF/RO_PSTA[20] , \REGF/RO_ACC[11] , \ADOSEL/n4120 , \LBUS/lnsa_end , 
        ph_lblockh, \LBUS/*cell*3982/U201/CONTROL1 , \PDOSEL/n115 , 
        \CODEIF/n3853 , \LBUS/n1400 , \CONS/n708 , \LBUS/n1590 , \CONS/n698 , 
        \SADR/pgaddwxz[6] , \pgsadrh[3] , \REGF/RO_ACC[22] , 
        \CODEIF/pgctrinc[17] , \pk_idcx_h[19] , \LDCHK/n3299 , \LDCHK/n3309 , 
        \ALUSHT/pkaluout[6] , \REGF/RI_SRA12M[12] , \pk_s1ba_h[15] , 
        \REGF/n8166 , \ALUSHT/pkshtout[3] , \LBUS/PIOSEL_1_Q1249 , 
        \PDOSEL/n225 , ph_sprlth, \pk_indz_h[8] , ph_exstgb_h, \REGF/n8141 , 
        \stream3[22] , \pk_rread_h[1] , \ADOSEL/n4097 , \ADOSEL/n4107 , 
        \CODEIF/n4004 , \ALUIS/n3739 , \pk_sra2_h[11] , \SADR/pgaddwz[23] , 
        \SADR/segbase[15] , \pk_s5ba_h[6] , \CODEIF/n3874 , \PDOSEL/n132 , 
        \LBUS/n1427 , \pk_idcy_h[16] , ph_adrdec_h, \REGF/RI_SRDA[3] , 
        \pk_pcs1_h[13] , \pk_s01l_h[22] , \CODEIF/n3968 , \BLU/n1551 , 
        \CONS/n633 , \stream3[20] , \stream3[13] , \pk_spr_h[8] , 
        \SADR/pgaddwz[10] , \pk_s01l_h[11] , \pk_sefl_h[5] , pktrscendh, 
        \REGF/pk_idcw_h[25] , \LDCHK/n3232 , \pk_adb_h[9] , \MAIN/n3616 , 
        ph_sa2lt_h, \pk_idcw_h[21] , \REGF/RO_LPSAS2156[4] , \pkbludgh[1] , 
        \SADR/pgaddwxy[7] , \SADR/pgaddwxz[4] , \pgsadrh[27] , \pgsadrh[14] , 
        \pk_sbba_h[9] , \pk_stdat[4] , \pgld32[12] , \CONS/n524 , \MAIN/n3631 , 
        \pk_s89l_h[24] , \pk_s89l_h[17] , \pk_idcw_h[12] , phatchkh, 
        \pk_s1ba_h[17] , \pk_s8ba_h[11] , \stream4[52] , \BLU/n1576 , 
        \pgld32[21] , \CONS/n614 , \LBUS/n1420 , \CONS/n728 , 
        \REGF/RI_SRA12M[23] , \REGF/RO_PSTA[22] , \CODEIF/n3873 , 
        \REGF/RO_ACC[13] , \PDOSEL/n135 , \ADOSEL/n4090 , \ADOSEL/n4100 , 
        \CODEIF/n4003 , \ALUSHT/pkshtout[1] , \REGF/RI_SRA12M[10] , 
        \REGF/n8146 , \pgsadrh[1] , ph_bitsrch, \CONS/n588 , \REGF/RO_ACC[20] , 
        \ALUSHT/pkaluout[4] , \CODEIF/pgctrinc[15] , \pk_s0ba_h[8] , 
        \pk_s45l_h[9] , \REGF/n8161 , \REGF/pk_scba_h[18] , \MAIN/reg_enable , 
        po_raccl_h, \MAIN/dprw_tap1 , \pk_sra2_h[20] , \pk_sra2_h[13] , 
        \pk_s5ba_h[4] , \LBUS/n1597 , \LBUS/n1407 , \PDOSEL/n112 , 
        \CODEIF/n3854 , \CODEIF/pfctr415[18] , \stream3[8] , \pk_dpr_h[31] , 
        \pk_dpr_h[28] , \SADR/pgaddyz[21] , \SADR/pgaddyz[12] , 
        \pk_rread_h[3] , \ALUIS/n3719 , \ADOSEL/n4127 , \CODEIF/n4024 , 
        \ALUIS/n3689 , \pgaluinb[6] , \pk_adb_h[21] , \CODEIF/pgfpce_in , 
        ph_errtendh, \pk_adb_h[12] , \pgaluina[5] , \pk_s2ba_h[16] , wspr, 
        \pk_sabl_h[0] , \ADOSEL/n4149 , \pk_rwrit_h[55] , \REGF/n8218 , 
        \REGF/RO_ERRA[10] , \CONS/n746 , \pk_rread_h[35] , \SADR/pgaddxyz[3] , 
        \pk_sfba_h[2] , \pk_pcs1_h[7] , \ALUIS/n3750 , \stream2[19] , 
        \pk_s67l_h[18] , \REGF/RO_ERRA[23] , \pk_rwrit_h[66] , \REGF/n8128 , 
        \MAIN/astregw_tap2 , \CODEQ/nqueue1[14] , \pk_idcz_h[20] , 
        \SADR/pgaddxz[9] , n10733, \SADR/operand[20] , \SADR/operand[5] , 
        \pk_sra1_h[7] , \SADR/pgaddwx[9] , \REGF/RO_TRCO[25] , \REGF/n8184 , 
        po_oprtrs_h, ph_exe_ah, \CODEQ/nqueue1[27] , \SADR/sadr[17] , 
        \pk_sdba_h[10] , \pk_scdl_h[19] , \LDIS/n3152 , \BLU/n1518 , 
        \CODEIF/n3921 , \BLU/n1488 , \pk_s45l_h[17] , \pk_sefl_h[28] , 
        ph_atchkenh, \pk_psae_h[6] , \pk_idcx_h[3] , \pk_sefl_h[31] , 
        \pkdptout[29] , \CODEIF/n3906 , \pk_s4ba_h[3] , \pkdptout[30] , 
        \CODEIF/n3896 , \pk_scdl_h[9] , \REGF/RO_ACC[7] , \stream3[1] , 
        \pk_dpr_h[21] , \pk_dpr_h[12] , \pk_indz_h[17] , \SADR/sadr[24] , 
        \REGF/pk_scti_h[0] , \pgmuxout[31] , \pgmuxout[28] , \pk_s45l_h[24] , 
        \pgaluina[18] , \CODEQ/nqueue2[57] , \pk_scba_h[7] , 
        \REGF/RO_PCON[24] , \pk_rread_h[16] , \stream2[10] , \CONS/n576 , 
        \pk_s67l_h[11] , \LDCHK/n3247 , \pk_rwrit_h[45] , \REGF/RO_ERRA[19] , 
        \pk_saco_hh[29] , \pk_rread_h[25] , \BLU/n1524 , \CONS/n646 , 
        \REG_2/n517 , \pk_s67l_h[22] , \pk_saco_hh[30] , \pk_spr_h[1] , 
        \pk_trba_h[8] , \SADR/pgaddwx[0] , \SADR/pgaddwyz[7] , \pk_s23l_h[2] , 
        \pk_sabl_h[9] , \REGF/RI_PCOH[5] , \REGF/RO_PCON[17] , \pk_stdat[15] , 
        \LDIS/n3149 , \CONS/n661 , \BLU/n1493 , \BLU/n1503 , \REGF/RO_EACC[6] , 
        \ALUIS/n3677 , \pk_adb_h[31] , \pk_adb_h[28] , \CONS/n340 , 
        \CONS/n551 , \MAIN/*cell*4603/U10/CONTROL1 , \SAEXE/n421 , 
        \pk_s1ba_h[6] , \pk_scdl_h[0] , \LDCHK/n3260 , \SAEXE/ph_lber1_h , 
        \REGF/n8133 , \pkdptout[13] , po_dprtrs_h, \pgmuxout[21] , 
        \pk_s6ba_h[12] , \pk_s01l_h[5] , \pk_sefl_h[21] , \pk_sefl_h[12] , 
        \pgaluina[11] , \CODEQ/nqueue2[47] , \pgaluina[22] , \PDOSEL/n96 , 
        \pgbluext[16] , \LBUS/n1455 , \PDOSEL/n140 , \pk_scdl_h[23] , 
        \pk_scdl_h[10] , \pk_idcw_h[7] , \REGF/RI_DPR[7] , \REGF/n8203 , 
        \pkdptout[20] , \pgmuxout[12] , \LDIS/ldexcl[4] , \CODEIF/n3996 , 
        \ADOSEL/n4152 , \CODEQ/nqueue1[37] , \REGF/pk_indz_h[30] , 
        \REGF/pk_indz_h[29] , \REGF/n8224 , wonly1, \pgbluext[3] , 
        \CONS/SACO[16] , \REGF/n8084 , \REGF/n8114 , \SADR/m_fadrl[7] , 
        \pgsdprlh[17] , \REGF/RO_LLPSAS[13] , \ALUIS/n3692 , \ALUIS/n3702 , 
        \pk_saco_lh[6] , po_ldis_h, \stream4[42] , ph_wdsrdaselh, \pgld32[31] , 
        \pgld32[28] , \CONS/n684 , \PDOSEL/n109 , \BLU/n1476 , \CONS/n714 , 
        ph_obmselh, \SADR/pgaddxz[14] , po_arsel_h, \MAIN/decend_en , 
        \LDCHK/n3285 , \SADR/pgaddwz[19] , \pgregadrh[17] , \pk_s5ba_h[13] , 
        \pkbludgh[8] , \pk_sbba_h[0] , \REGF/pk_idcy_h[31] , 
        \REGF/pk_idcy_h[28] , \pk_s89l_h[6] , \pk_adb_h[0] , \CONS/n593 , 
        \SADR/pgaddwxy[21] , \SADR/pgaddwxy[12] , \SADR/lmtaddr[11] , 
        \pk_s01l_h[18] , \pk_sabl_h[27] , \pk_s67l_h[7] , \CODEIF/n4018 , 
        \ALUIS/n3725 , \pk_sabl_h[14] , \REGF/RI_SPR[2] , \CODEIF/n3868 , 
        \CODEIF/pfctr415[4] , \CONS/n733 , \REGF/pk_idcx_h[25] , \LDIS/n3127 , 
        pk_bitdatah, \CODEIF/n3954 , \SADR/operand[13] , \stream3[30] , 
        \PDOSEL/n182 , \stream3[29] , \pk_indz_h[3] , \pk_s45l_h[0] , 
        \CODEIF/pfctr415[11] , ph_pdlen_h, \pk_sra2_h[30] , \pk_sra2_h[29] , 
        \REGF/n8061 , \pk_s0ba_h[1] , \REGF/RI_SRA12M[19] , \REGF/RO_PSTA[18] , 
        ph_ltwt_h, \ALUSHT/pkshtout[8] , \SADR/operand[1] , \pk_indz_h[20] , 
        \pgsadrh[8] , \pk_idcx_h[12] , \LBUS/n1610 , \CONS/n518 , 
        \SADR/sadr[13] , \pk_s4ba_h[7] , \pk_scba_h[15] , \pk_s23l_h[24] , 
        \pgsdprlh[5] , \REGF/RO_ACC[29] , \pk_s23l_h[17] , \REGF/RO_ACC[30] , 
        \pk_idcx_h[21] , \CODEIF/n3973 , \MAIN/POL_STH , \CONS/n628 , 
        \pk_idcy_h[5] , \REGF/RO_ACC[3] , \CODEIF/wprotect0 , \LDIS/ldexcl[9] , 
        \CODEIF/n3946 , \pk_s01l_h[8] , \pk_s45l_h[13] , \LDIS/n3135 , 
        \pk_indz_h[13] , \pk_sdba_h[14] , \pk_psae_h[2] , \pk_idcx_h[7] , 
        \pk_s45l_h[20] , \CODEQ/nqueue2[53] , \SADR/sadr[20] , \REGF/n8073 , 
        \REGF/pk_scti_h[4] , \pgbluext[31] , \pgbluext[28] , \stream3[24] , 
        \stream3[17] , \pk_sra1_h[3] , \REGF/pk_indz_h[24] , \REGF/n8054 , 
        mem_cnfg_h, \LBUS/n1602 , ronly2, \CODEIF/n3961 , word32odtrh, 
        \CODEQ/nqueue1[10] , \BLU/n1558 , ph_sprtrs_h, \SADR/pgaddyz[16] , 
        \SADR/pgaddxyz[7] , \pk_sfba_h[6] , \CODEQ/nqueue1[23] , 
        \REGF/RI_PCOH[8] , \pk_rwrit_h[51] , \pk_rwrit_h[48] , \pk_pcs1_h[3] , 
        \ALUIS/n3680 , \ALUIS/n3710 , \REGF/RO_ERRA[14] , \pk_rread_h[31] , 
        \pk_rread_h[28] , \CONS/n696 , \CONS/n706 , \REGF/n_2734 , 
        \REGF/RO_ERRA[27] , \BLU/n1464 , \REGF/RO_PCON[30] , \LDCHK/n3297 , 
        \LDCHK/n3307 , \REGF/RO_PCON[29] , \REGF/n8168 , \pk_rwrit_h[62] , 
        \pgaluina[1] , \pk_adb_h[25] , \pgaluinb[2] , \CONS/n581 , 
        \pk_s2ba_h[12] , \pk_sabl_h[4] , \pk_stdat[18] , po_lwdsrc_h, 
        \ADOSEL/n4109 , \ADOSEL/n4099 , accbsel, \ALUIS/n3737 , \LBUS/n1429 , 
        \CONS/n721 , \pk_adb_h[16] , \CODEIF/fadren , \pk_rread_h[7] , 
        \REGF/n8121 , \pk_sra2_h[17] , \pk_trba_h[5] , \SADR/pgaddxz[19] , 
        \SADR/pgaddwxy[3] , \pk_s5ba_h[0] , \pk_s8ba_h[15] , \REGF/n8211 , 
        \CODEIF/n3984 , \REGF/RI_SRA12M[27] , \LBUS/n1447 , \PDOSEL/n152 , 
        \REGF/pk_idcx_h[31] , \REGF/pk_idcx_h[28] , \pk_idcy_h[8] , 
        \ADOSEL/n4140 , \CODEIF/n4043 , \REGF/RO_ACC[17] , \REGF/n8236 , 
        \pgsdprlh[8] , \LBUS/n1460 , \SADR/pgaddwxz[0] , \pgsadrh[5] , 
        \pk_s23l_h[30] , \pk_s23l_h[29] , \CODEIF/pgctrinc[11] , 
        \REGF/RO_ACC[24] , \ALUSHT/pkaluout[0] , ph_btsrdaselh, \REGF/n8106 , 
        \pgsadrh[10] , \pk_s1ba_h[13] , \REGF/RI_SRA12M[14] , \REGF/n8096 , 
        \ALUSHT/pkshtout[5] , \pk_s89l_h[20] , \pk_stdat[0] , \pgld32[16] , 
        \CONS/n564 , \SAEXE/n414 , \REGF/pk_idcy_h[25] , \pkbludgh[5] , 
        \LDCHK/n3255 , \REGF/RO_LPSAS2156[0] , \pgsadrh[23] , \pk_s89l_h[13] , 
        \stream4[56] , rmw11, \CONS/n654 , \pgld32[25] , \BLU/n1536 , 
        \pk_s01l_h[26] , \pk_idcw_h[16] , \MAIN/cstregw_tap1 , \CONS/n673 , 
        \pk_sabl_h[19] , \BLU/n1481 , \BLU/n1511 , \RSTGN/CRST_1H , 
        \SADR/pgaddwz[14] , \SADR/segbase[11] , \REGF/RI_SRDA[7] , 
        \CODEIF/pfctr415[9] , \CODEIF/n3928 , \pk_pcs1_h[17] , \pk_idcy_h[12] , 
        \ALUIS/n3665 , \REGF/pk_exco_h[2] , \pk_s01l_h[15] , \pk_sefl_h[1] , 
        \pk_idcy_h[21] , \LDCHK/n3272 , \CONS/n543 , \SADR/operand[24] , 
        \SADR/pgaddwxz[9] , \pk_scba_h[11] , \pk_s23l_h[20] , \pgsdprlh[1] , 
        ph_ldaoutenh4, \CODEIF/pgctrinc[18] , \LDCHK/n3269 , \SAEXE/n428 , 
        \pk_idcx_h[16] , \ALUSHT/pkaluout[9] , \CONS/n349 , \CONS/n558 , 
        \pk_s5ba_h[9] , \pk_s23l_h[13] , \pk_idcy_h[1] , \REGF/n8196 , 
        \REG_2/ncnt1[0] , \CODEIF/n3933 , \CONS/n668 , \ALUIS/n3659 , 
        \LDIS/n3140 , \CODEIF/pfctr415[15] , \stream3[34] , \CODEIF/n3884 , 
        \SADR/operand[17] , \pk_s0ba_h[5] , \CODEIF/n3914 , ph_lbslock_h, 
        \REGF/pk_s8ba_h[18] , \SADR/operand[8] , \pk_spr_h[5] , 
        \SADR/pgaddxz[23] , \SADR/pgaddwxy[16] , \pk_indz_h[7] , 
        \pgregadrh[13] , \pk_s45l_h[4] , po_shelter_h2, \pk_sabl_h[23] , 
        \pk_s89l_h[2] , \pk_sefl_h[8] , \pk_adb_h[4] , \REGF/pk_idcw_h[31] , 
        \REGF/pk_idcw_h[28] , \pgregadrh[20] , \SADR/lmtaddr[15] , 
        \pk_s67l_h[3] , \pk_sabl_h[10] , \REGF/RI_SPR[6] , 
        \CODEIF/pfctr415[0] , \BLU/n1581 , \pk_saco_lh[2] , \stream4[46] , 
        po_cmfsel_h, \PDOSEL/n149 , \pgsadrh[19] , \pk_sbba_h[4] , 
        \pgsdprlh[13] , \ALUIS/n3742 , \pk_s89l_h[30] , \pk_s89l_h[29] , 
        \pk_stdat[9] , \SADR/pgaddwx[4] , \SADR/pgaddxz[10] , \pk_s5ba_h[17] , 
        \pgsdprlh[20] , \pk_scdl_h[14] , \REGF/RO_LPSAS2156[9] , 
        \pk_idcw_h[3] , \REGF/RO_DDCS[25] , \pgbluext[7] , \CODEIF/n3861 , 
        \PDOSEL/n127 , \CONS/SACO[12] , \LBUS/n1432 , \REGF/RI_DPR[3] , 
        pk_bacch, \ADOSEL/n4112 , \CODEIF/n4011 , \CODEQ/nqueue1[33] , 
        \pk_s1ba_h[2] , \pk_s45l_h[30] , \pk_s45l_h[29] , \pk_scdl_h[27] , 
        \REGF/n8154 , \CODEQ/nqueue1[19] , \pk_sefl_h[16] , \pgmuxout[25] , 
        \pgaluina[15] , \CODEQ/nqueue2[43] , \REGF/n8173 , \pkdptout[17] , 
        \stream3[5] , \pk_dpr_h[16] , \SADR/pgaddwyz[3] , \pk_s6ba_h[16] , 
        \pk_scdl_h[4] , \pkdptout[24] , \REGF/n8243 , \CODEIF/n3846 , 
        \pgmuxout[16] , \LDIS/ldexcl[0] , \PDOSEL/n100 , \pk_s01l_h[1] , 
        \pgaluina[26] , \LBUS/n1415 , \pk_s23l_h[6] , \pk_sefl_h[25] , 
        pgadrovfh, \ADOSEL/n4135 , \CODEIF/n4036 , \pk_stdat[11] , 
        \REGF/RO_EACC[2] , \pgaluina[8] , \CONS/n621 , \BLU/n1543 , pk_pcsee_h, 
        \pk_scba_h[3] , \pk_s67l_h[15] , \CONS/n300 , ph_dec_bh, 
        \REGF/RO_PCON[20] , \pk_rread_h[12] , \REGF/n8068 , \MAIN/n3623 , 
        \stream2[14] , \REGF/RI_PCOH[1] , \CONS/n536 , \REGF/RO_PCON[13] , 
        \SADR/pgaddwy[22] , \SADR/pgaddwy[11] , \SADR/pgaddxz[4] , 
        \pk_s67l_h[26] , \pk_rwrit_h[41] , pk_sased_h, \CONS/n606 , 
        \pk_rread_h[38] , \pk_rread_h[21] , \stream2[27] , \pk_rwrit_h[58] , 
        \BLU/n1564 , \pk_pdo_h[4] , phlmterr_h, \PDOSEL/n108 , \BLU/n1477 , 
        \CONS/n685 , \CONS/n715 , \stream4[23] , step4_cf, \ALUIS/n3693 , 
        \ALUIS/n3703 , \SADR/pgaddxy[7] , \pk_saba_h[13] , \stream4[6] , 
        \pgldi[27] , \ALUSHT/pkshtout[31] , \ALUSHT/pkshtout[28] , 
        \REGF/RI_PCOL[1] , \stream4[10] , \LBUS/flag_tr2 , \REGF/RI_TBAI[9] , 
        \pgldi[14] , \SADR/pgovfxz , \pk_seba_h[5] , \LDCHK/n3284 , 
        \CONS/n592 , \ph_pdis_h[3] , \pk_spr_h[31] , \pk_spr_h[28] , 
        \pk_sra1_h[19] , \SADR/pgaddwy[9] , \SADR/pgovfwxyz , 
        \REGF/RI_TBAI[16] , \REGF/RO_SRDA[1] , \pk_pc_h[7] , \CODEIF/n3869 , 
        \CODEQ/nqueue1[7] , \CONS/n732 , \CODEIF/n4019 , \ALUIS/n3724 , 
        \CODEQ/nqueue2[4] , \pk_pc_h[11] , \REGF/RI_DPR[23] , \stream3[51] , 
        \stream3[48] , \pgld16[13] , \MAIN/sprw_tap1 , \pk_s9ba_h[1] , 
        \REGF/RI_SRDA[30] , \REGF/RI_SRDA[29] , \LDIS/n3126 , \CODEIF/n3955 , 
        \PDOSEL/n183 , \REGF/RI_DPR[10] , \LDCHK/pglpinff[3] , 
        \SADR/pgaddwxyz[21] , \pk_indw_h[4] , \pk_indx_h[10] , \pk_indx_h[9] , 
        \SADR/segbase[6] , \REGF/n8060 , \REGF/RI_ACC[22] , \pk_s7ba_h[4] , 
        \pk_s2ba_h[8] , \pk_s7ba_h[15] , \REGF/RO_EACC[26] , \REGF/RI_STAT[3] , 
        \UPIF/ph_accessenh , \LBUS/n1611 , \CONS/n519 , \CONS/n298 , 
        \REGF/RI_ACC[11] , \CODEIF/wprotect1 , \REGF/RO_EACC[15] , \CONS/n629 , 
        \REGF/RI_SPR[22] , \CODEIF/n3972 , \LDCHK/n3246 , \LBUS/ilt[4] , 
        \SADR/pgaddwxyz[4] , \CONS/n577 , \pgldi[6] , \pk_spr_h[21] , 
        \pk_spr_h[12] , \pk_dpr_h[0] , \pk_trba_h[31] , \pk_trba_h[28] , 
        \pk_rwrit_h[17] , \ALUIS/n3651 , \SADR/pgaddwxyz[12] , \pk_indx_h[23] , 
        \REGF/RI_SPR[11] , \SADR/lmtaddr[3] , \pk_rread_h[44] , 
        \pk_rwrit_h[24] , \CODEIF/pgctrinc[5] , \pkbludgh[14] , 
        \LBUS/*cell*3982/U158/Z_0 , \BLU/n1525 , \pk_trba_h[21] , 
        \SADR/pgaddwyz[15] , \pk_s4ba_h[14] , \REGF/RI_PCOH[18] , 
        \REGF/pk_indx_h[27] , \CONS/n647 , \stream1[18] , \ALUIS/n3676 , 
        \pk_sdba_h[2] , \REGF/RO_PSASL[1] , \CODEIF/pfctr[10] , 
        \MAIN/*cell*4603/U14/CONTROL1 , \pgld32[8] , \BLU/n1492 , \BLU/n1502 , 
        \REGF/RO_PCON[0] , \LDIS/n3148 , \CONS/n660 , \pk_saco_lh[14] , 
        \LDCHK/n3261 , \pk_ada_h[5] , \SAEXE/n420 , ph_word16_h, \CONS/n550 , 
        \CONS/n341 , \pk_indw_h[19] , \pk_indy_h[6] , \pk_ada_h[18] , 
        \REGF/n8132 , \pk_s8ba_h[6] , \pk_sbba_h[12] , \REGF/RI_PCOL[30] , 
        \REGF/RI_EACC[30] , \REGF/RI_EACC[29] , \CODEQ/nqueue2[26] , 
        \REGF/n8202 , \CODEIF/pfctr[6] , \ALUSHT/pkaluout[26] , \CODEIF/n3997 , 
        \LBUS/n1454 , \CODEQ/nqueue2[15] , \PDOSEL/n97 , \PDOSEL/n141 , 
        \REGF/RI_PCOL[29] , \REGF/RO_SRDA[26] , \REGF/RO_LLPSAS[7] , 
        ph_stage_ah, \ALUSHT/pkaluout[15] , \REGF/n8225 , \pk_s6ba_h[3] , 
        \pk_idcz_h[0] , \ADOSEL/n4153 , \pgaluinb[19] , \CODEQ/nqueue1[56] , 
        \pk_saba_h[7] , \REGF/RI_PCOH[22] , \REGF/RO_SRDA[15] , \REGF/n8115 , 
        \REGF/RO_PPCN[10] , \REGF/n8085 , \pkdptout[0] , \REGF/RO_PCON[9] , 
        \REGF/RI_PCOH[11] , \REGF/RI_SRA12M[5] , \pk_ada_h[11] , \stream1[22] , 
        \ph_cpudout[4] , \CONS/SACO[3] , \stream1[11] , \ADOSEL/n4148 , 
        \pgld32[1] , \pk_sfba_h[16] , \REGF/RO_PSASL[8] , \REGF/RI_EACC[4] , 
        \pk_ada_h[22] , \REGF/RI_SPR[18] , \ALUIS/n3751 , \ph_cpudout[15] , 
        \pk_dpr_h[9] , \pk_pdo_h[17] , \pk_rwrit_h[34] , \REGF/n8219 , 
        \CONS/n747 , \pk_trba_h[12] , ph_stregwt_h, \pk_rread_h[54] , 
        \REG_2/RETCNT[4] , \pk_indx_h[19] , \ph_cpudout[26] , \pk_pdo_h[24] , 
        \SADR/pgaddwx[21] , \SADR/pgaddwx[12] , \pk_indw_h[23] , \REGF/n8185 , 
        \REGF/n8129 , \phshtd[5] , \pk_indw_h[10] , \pkdptout[9] , 
        \pgaluinb[23] , \LDIS/n3153 , \BLU/n1489 , \pk_indy_h[14] , 
        \pk_s3ba_h[6] , \CODEIF/n3920 , \BLU/n1519 , \pk_idcz_h[9] , 
        \CODEQ/nqueue1[46] , \pgaluinb[10] , \pk_s0ba_h[10] , 
        \REGF/RI_EACC[13] , \SADR/pgaddyz[7] , \SADR/pgaddxyz[15] , 
        \ph_segset_h[6] , \REGF/RI_PCOL[20] , \CODEIF/n3897 , \CODEIF/n3907 , 
        \pk_s9ba_h[16] , \pgld16[7] , \REG_2/ph_retcnt_h[6] , 
        \REGF/pk_indw_h[27] , \SADR/pgaddxy[15] , \REGF/RI_PCOL[13] , 
        \REGF/RI_EACC[20] , \CODEQ/nqueue2[36] , \CODEIF/frpend_in , 
        \stream2[1] , \CODEIF/n3969 , \LDIS/ldexcl[15] , \REGF/RO_SRDA[8] , 
        oebacc, \CONS/n632 , \BLU/n1550 , \REGF/RO_PPCN[4] , \stream1[2] , 
        \SAEXE/sa_start1 , \MAIN/n3617 , \pk_dpr_h[4] , \pk_sra1_h[23] , 
        \pk_sra1_h[10] , \pk_sra2_h[2] , \SADR/pgaddwy[18] , 
        \SADR/pgaddwxz[13] , \ph_segset_h[24] , \pk_pcs2_h[10] , 
        \pk_idcz_h[15] , \LDCHK/n3233 , \stream4[19] , \ALUSHT/pkshtout[21] , 
        \CONS/n525 , \MAIN/n3630 , \pk_s3ba_h[11] , \ph_segset_h[17] , 
        \REGF/RI_PCOL[8] , \REGF/RI_TBAI[0] , \REGF/RO_EST1[0] , \stream4[33] , 
        \BLU/n1577 , \ALUSHT/pkshtout[12] , \pk_rwrit_h[2] , \CONS/n615 , 
        \pk_pcs2_h[2] , \SADR/pgaddwxz[20] , \pk_s2ba_h[1] , \REGF/RI_ACC[5] , 
        \REGF/RO_ERRA[7] , \ADOSEL/n4101 , \pgmuxout[4] , \ADOSEL/n4091 , 
        \REGF/RI_ACC[18] , \CODEIF/n4002 , \SADR/pgaddwy[0] , \pk_indx_h[0] , 
        \pk_seba_h[17] , \CODEIF/n3872 , \LDCHK/lpex[3] , \LBUS/n1421 , 
        \CONS/n729 , \PDOSEL/n134 , pk_pcovf_h, \REGF/RI_DPR[19] , 
        \REGF/n8147 , srctype2, \CONS/n589 , \SADR/pgaddwz[3] , 
        \REGF/RI_SRDA[13] , \REGF/pk_s7ba_h[18] , \REGF/n8160 , \PDOSEL/n223 , 
        \stream3[58] , \LDIS/ldexch[17] , \SADR/pgaddwyz[22] , 
        \SADR/pgaddxyz[18] , \pk_indy_h[2] , \SADR/m_fadrl[15] , 
        \REGF/RI_SRDA[20] , \pk_pc_h[18] , \stream3[41] , \CODEIF/n4025 , 
        \ALUIS/n3688 , \ALUIS/n3718 , \ADOSEL/n4126 , \pk_s6ba_h[7] , 
        \pk_s9ba_h[8] , \pgregadrh[3] , \LDIS/ldexch[24] , \LBUS/n1406 , 
        \LBUS/n1596 , \REGF/RO_SRDA[22] , \pk_idcz_h[4] , \ADOSEL/n4113 , 
        \CODEIF/n3855 , \PDOSEL/n113 , \CODEIF/n4010 , \CODEQ/nqueue1[52] , 
        \CODEIF/n3860 , \PDOSEL/n126 , \REGF/RO_SRDA[11] , \REGF/RO_PPCN[14] , 
        ph_sastlth, \LBUS/n1433 , \REGF/n8155 , \pkdptout[4] , 
        \CODEIF/pfctr[2] , \poalufnc[2] , \ALUSHT/pkaluout[22] , \LBUS/MMBSEL , 
        \CODEQ/nqueue2[22] , \REGF/n8172 , \ADOSEL/n4134 , \pk_indy_h[19] , 
        \pk_s8ba_h[2] , \CODEIF/n4037 , \ALUSHT/pkaluout[11] , \pk_sbba_h[16] , 
        ph_lmterr_h, \REGF/n8242 , \CODEIF/n3847 , \LBUS/n1395 , \PDOSEL/n101 , 
        \LBUS/n1414 , \CODEQ/nqueue2[11] , \CONS/n620 , \BLU/n1542 , 
        \SADR/pgaddwyz[11] , \pk_s4ba_h[10] , \pk_sati_h[0] , 
        \REGF/RI_EACC[9] , \REGF/RI_SRA12M[8] , \pk_saco_lh[23] , 
        \CODEIF/pfctr[14] , \SADR/pgaddwxyz[0] , \pk_sdba_h[6] , 
        \pk_saco_lh[10] , \pk_ada_h[1] , \SAEXE/exec_end1 , \ph_cpudout[9] , 
        \pk_rwrit_h[13] , \REGF/RO_PCON[4] , \REGF/n8069 , ph_lpdilth, 
        \MAIN/n3622 , \pk_indx_h[14] , \pgldi[2] , \pk_pdo_h[30] , \CONS/n537 , 
        \pk_pdo_h[29] , \LBUS/ilt[0] , pk_pexe01_h, \REGF/RI_SPR[26] , 
        \CODEIF/wpfcinc , \SADR/pgaddwxyz[16] , \CONS/n607 , \pk_indw_h[0] , 
        \SADR/m_fadrl[18] , \SADR/segbase[2] , \SADR/lmtaddr[7] , 
        \pk_rread_h[59] , \pk_rread_h[40] , \pk_s7ba_h[11] , \pk_rwrit_h[39] , 
        \pk_rwrit_h[20] , \BLU/n1565 , \CODEIF/pgctrinc[1] , \pkbludgh[10] , 
        \REGF/RI_SPR[15] , \CONS/n348 , \ph_cpudout[18] , \CONS/n559 , 
        \pk_s7ba_h[0] , \REGF/RO_EACC[22] , \REGF/n8197 , \pk_s9ba_h[5] , 
        \REGF/RO_EACC[11] , \REGF/RI_ACC[26] , \LDCHK/n3268 , \SAEXE/n429 , 
        \CODEIF/n3932 , \REGF/RI_ACC[15] , \LDIS/n3141 , \CONS/n669 , 
        \REGF/RI_ACC[8] , \pgmuxout[9] , \CODEIF/n3885 , \CODEIF/n3915 , 
        \LDIS/ldexch[30] , \LDIS/ldexch[29] , \pk_pc_h[15] , \REGF/RI_DPR[27] , 
        \ALUIS/n3658 , \stream3[55] , \pk_idcz_h[18] , \REGF/RI_DPR[14] , 
        \SADR/m_fadrh[30] , \pk_seba_h[1] , \REGF/RI_TBAI[21] , 
        \REGF/pk_s3ba_h[18] , \ph_pdis_h[7] , \REGF/RO_SRDA[5] , 
        \REGF/RO_PPCN[9] , \pk_pc_h[3] , \CODEQ/nqueue1[3] , 
        \CODEQ/nqueue2[0] , \SADR/m_fadrh[29] , \pk_sra1_h[14] , 
        \SADR/pgaddwy[15] , \SADR/pgaddxy[18] , \SADR/pgaddxy[3] , 
        \REGF/RI_TBAI[12] , \BLU/n1580 , \pgldi[23] , \SADR/pgaddwz[7] , 
        \SADR/pgaddxz[0] , \ALUIS/n3743 , \pk_pdo_h[0] , \stream4[27] , 
        \PDOSEL/n148 , \SADR/m_fadrl[22] , \pk_saba_h[17] , \ph_segset_h[30] , 
        \pgldi[10] , \MAIN/single_read , \REGF/RI_PCOL[5] , \ph_segset_h[29] , 
        \stream4[2] , \stream4[14] , \REGF/RI_SRDA[17] , \pk_indw_h[9] , 
        \REGF/n8120 , \pk_sra2_h[6] , \SADR/pgaddwy[4] , \SADR/m_fadrl[11] , 
        \SADR/intbitno[2] , \REGF/n8210 , \CODEIF/n3985 , lbus_start, 
        \PDOSEL/n153 , \pgregadrh[7] , \REGF/RI_SRDA[24] , \LDIS/ldexch[20] , 
        \LBUS/n1446 , \REGF/RO_EACC[18] , \stream3[45] , \REGF/n8237 , 
        \SADR/pgaddwxz[17] , \pk_indx_h[4] , \pk_s2ba_h[5] , \CODEIF/n4042 , 
        \LBUS/n1461 , \REGF/RO_ERRA[3] , \ADOSEL/n4141 , \pgmuxout[0] , 
        ph_izco_h, \REGF/RI_ACC[1] , \REGF/n8097 , \REGF/n8107 , 
        \pk_s7ba_h[9] , \pk_seba_h[13] , \REGF/RI_TBAI[4] , \pgldi[19] , 
        \LDCHK/n3254 , \SAEXE/n415 , \REGF/RO_EST1[4] , \pgbitnoh[1] , 
        \pk_s3ba_h[15] , \MAIN/astregw_inhibith , \ALUSHT/pkshtout[25] , 
        \CONS/n565 , \ph_segset_h[20] , \ph_segset_h[13] , \pk_rwrit_h[6] , 
        \pk_pcs2_h[6] , st_cfctl, \REGF/pk_idcz_h[26] , \ALUIS/n3643 , 
        \CONS/n655 , \pk_pdo_h[9] , \stream4[37] , \ALUSHT/pkshtout[16] , 
        \BLU/n1537 , n10732, \pk_idcz_h[22] , \ALUIS/n3664 , \MAIN/ph_rmw1h , 
        ph_ex2regwt_h, \CODEQ/nqueue2[9] , \CONS/n672 , \SADR/pgaddxy[11] , 
        \pk_pcs2_h[14] , \pk_idcz_h[11] , \CODEIF/n3929 , \LDIS/ldexcl[11] , 
        \BLU/n1480 , \BLU/n1510 , \LDCHK/n3273 , n10735, \RSTGN/WRST_1H , 
        \pk_spr_h[16] , \SADR/pgaddwx[16] , \SADR/pgaddxy[22] , \pk_seba_h[8] , 
        step1_cf, \SADR/pgaddyz[3] , \SADR/pgaddxyz[11] , \ph_segset_h[2] , 
        \REGF/RO_PPCN[0] , baccsel, ph_mmbselh, \pgld16[3] , \CONS/n542 , 
        \ALUSHT/pkaluout[18] , \REGF/RI_PCOL[24] , \CODEIF/n3947 , 
        \SADR/pgaddxyz[22] , \pk_indy_h[10] , \pk_s0ba_h[14] , \LDIS/n3134 , 
        \REGF/RI_EACC[17] , \MAIN/st_decctl , \REGF/RI_PCOL[17] , 
        \CODEQ/nqueue2[18] , \pk_indw_h[14] , \pk_indy_h[23] , 
        \REGF/RI_EACC[24] , sequencial2, \CODEQ/nqueue2[32] , \pk_s3ba_h[2] , 
        \pk_s9ba_h[12] , \REGF/n8072 , \REGF/RO_SRDA[18] , 
        \REGF/pk_indy_h[27] , \pgaluinb[27] , \REG_2/ph_retcnt_h[2] , 
        \LBUS/n1603 , \REGF/n8055 , \phshtd[1] , \pgaluinb[14] , 
        \CODEQ/nqueue1[42] , \CODEIF/n3960 , \pk_rread_h[50] , exetype1, 
        \BLU/n1559 , \LDIS/n3113 , \pk_rread_h[49] , \pk_pdo_h[13] , 
        \CONS/n697 , \CONS/n707 , \pk_rwrit_h[30] , \pk_rwrit_h[29] , 
        \BLU/n1465 , \pk_trba_h[16] , \SADR/pgaddwxyz[9] , 
        \CODEIF/pgctrinc[8] , \ALUIS/n3681 , \ALUIS/n3711 , \ph_cpudout[11] , 
        rrmw2, \pk_pdo_h[20] , \REGF/n8169 , \pk_rread_h[63] , \LDCHK/n3296 , 
        \ph_cpudout[22] , \LDCHK/n3306 , \SADR/pgaddwx[14] , 
        \SADR/pgaddwyz[18] , \REGF/RI_SRA12M[1] , \REG_2/RETCNT[0] , 
        \pk_indy_h[12] , \pk_s0ba_h[16] , \pk_saba_h[3] , \pk_sfba_h[12] , 
        \REGF/RI_PCOH[26] , \pk_saco_lh[19] , \pk_ada_h[15] , \pk_ada_h[8] , 
        \stream1[26] , \CONS/SACO[7] , \CONS/n580 , \ph_cpudout[0] , 
        \LBUS/n1428 , \CONS/n720 , \pk_ada_h[26] , ph_lockh, 
        \REGF/RI_PCOH[15] , \REGF/RI_EACC[0] , \ADOSEL/n4098 , \pgld32[5] , 
        \stream1[15] , \ADOSEL/n4108 , \ALUIS/n3736 , \REGF/RI_EACC[15] , 
        \CODEIF/n3967 , \LDIS/n3114 , \SADR/pgaddyz[1] , \SADR/pgaddxyz[13] , 
        \pk_s8ba_h[9] , \REG_2/ncnt3[1] , \REGF/RI_PCOL[26] , 
        \SADR/pgaddxyz[20] , \pk_indy_h[21] , \pk_indy_h[9] , \pk_s9ba_h[10] , 
        \ph_segset_h[0] , \pgld16[1] , \LBUS/OBMSEL , \REGF/n8052 , allfbsel, 
        \MAIN/n3619 , \REG_2/ph_retcnt_h[0] , \REGF/RI_EACC[26] , \LBUS/n1604 , 
        \CODEQ/nqueue2[30] , \CODEIF/pgfpoe_in , \ALUSHT/pkaluout[30] , 
        \CODEQ/nqueue2[29] , \ALUSHT/pkaluout[29] , \REGF/RI_PCOL[15] , 
        \REGF/pk_indy_h[25] , \REGF/n8075 , immbsel, \CODEIF/pfctr[9] , 
        \phshtd[3] , \CODEIF/fm_config[1] , \pgaluinb[25] , \pk_spr_h[14] , 
        \pk_indw_h[16] , \REGF/RO_LLPSAS[8] , \LDIS/n3133 , \pk_s3ba_h[0] , 
        \BLU/n1579 , ph_lbe3_h, \REGF/RO_SRDA[30] , \REGF/RO_SRDA[29] , 
        \CODEIF/n3940 , pk_rgbit_h, \pgaluinb[16] , \CODEQ/nqueue1[59] , 
        \CODEQ/nqueue1[40] , \ALUIS/n3731 , \ph_cpudout[13] , \pk_trba_h[14] , 
        ph_wrdsrc_h, \pk_rread_h[52] , \pk_pdo_h[11] , \pk_rwrit_h[32] , 
        \CONS/n727 , \REG_2/RETCNT[2] , \ph_cpudout[20] , \SADR/pgaddwy[6] , 
        \pk_saba_h[1] , \pgldi[9] , \pk_rread_h[61] , \REGF/RI_PCOH[24] , 
        \pk_rwrit_h[18] , \pk_pdo_h[22] , \CONS/n587 , \REGF/n8149 , 
        \REGF/RI_PCOH[17] , \REGF/RI_SRA12M[3] , \pk_ada_h[17] , \LDCHK/n3291 , 
        \LDCHK/n3301 , \ph_cpudout[2] , \CONS/SACO[5] , \ALUIS/n3686 , 
        \ALUIS/n3716 , \REGF/pk_indx_h[28] , \REGF/pk_indx_h[31] , 
        \REGF/RI_EACC[2] , \ADOSEL/n4128 , \pgld32[7] , \pk_sfba_h[10] , 
        \pk_ada_h[24] , \LBUS/n1408 , \CONS/n700 , \LBUS/n1598 , \CONS/n690 , 
        \pk_sra1_h[16] , \pk_sra2_h[4] , \SADR/pgaddwz[5] , \REGF/RI_SRDA[15] , 
        \REGF/n8090 , \REGF/n8100 , \SADR/m_fadrl[20] , \SADR/m_fadrl[13] , 
        saenabl1, \stream3[47] , \ADOSEL/n4146 , \LDIS/ldexch[22] , 
        \SADR/intbitno[0] , \pgregadrh[5] , \REGF/RI_SRDA[26] , \LBUS/EXTSEL , 
        \pk_s2ba_h[7] , \REGF/pk_stat_h[16] , \REGF/RI_ACC[3] , \REGF/n8230 , 
        \REGF/RO_ERRA[1] , \pgmuxout[2] , pol_status, \CONS/n749 , 
        \SADR/pgaddwxz[15] , \pk_indx_h[6] , \SADR/segbase[9] , \REGF/n8217 , 
        \CODEIF/n3982 , \LBUS/n1441 , \PDOSEL/n82 , \PDOSEL/n154 , 
        \pk_seba_h[11] , \pgbitnoh[3] , \REGF/RO_EACC[30] , \REGF/RO_EACC[29] , 
        \REGF/n8127 , \pk_s3ba_h[17] , \ph_segset_h[22] , \CONS/n545 , 
        \REGF/RO_EST2[5] , \stream4[9] , all0asel, \ALUSHT/pkshtout[27] , 
        \REGF/RI_TBAI[6] , \REGF/RO_EST1[6] , \LDCHK/n3274 , \BLU/n1487 , 
        pgfbadrsel, \stream4[35] , \ALUSHT/pkshtout[14] , \BLU/n1517 , 
        \CONS/n675 , \SADR/pgaddxy[13] , \SADR/pgaddxy[8] , \ph_segset_h[11] , 
        \pk_rwrit_h[4] , \pk_pcs2_h[4] , pr_write_h, \ALUIS/n3663 , 
        \REGF/pk_idcz_h[24] , \REGF/RI_TBAI[19] , \pgldi[31] , \pgldi[28] , 
        \CODEIF/n3899 , \CODEIF/n3909 , \LDIS/ldexcl[13] , \pk_pc_h[8] , 
        \CODEQ/nqueue1[8] , \BLU/n1530 , \CONS/n652 , \SADR/pgaddxy[20] , 
        \REGF/RO_PPCN[2] , \REGF/pk_saba_h[18] , \LBUS/nlt[0] , \CONS/n562 , 
        \SADR/pgovfwz , \pk_indw_h[2] , \SADR/segbase[0] , \pk_pcs2_h[16] , 
        \pk_idcz_h[13] , \LDCHK/n3253 , \SAEXE/n412 , \REGF/RI_ACC[24] , 
        \pk_s7ba_h[13] , \pk_s7ba_h[2] , \LDCHK/n3248 , \REGF/RO_EACC[20] , 
        \REGF/RI_STAT[5] , ebaccsel, \pk_s9ba_h[7] , \REGF/RO_ERRA[8] , 
        \REGF/RI_ACC[17] , \LBUS/*cell*3982/U188/CONTROL1 , \CONS/n579 , 
        \pk_pc_h[17] , \REGF/RO_EACC[13] , \LDIS/n3161 , \CONS/n649 , 
        \REGF/RI_DPR[25] , \stream3[57] , \CODEIF/n3882 , \CODEIF/n3912 , 
        \MAIN/EXCEP_EXT , \pgld16[15] , \ALUIS/n3678 , \CODEIF/n3935 , 
        \LDIS/n3146 , \REGF/RI_DPR[16] , ph_ldaoutenh2, \pk_seba_h[3] , 
        ph_tbllt_h, \REGF/n8190 , \LDIS/ldexch[18] , \ALUSHT/aluovf , 
        \REGF/RI_TBAI[23] , \ph_pdis_h[5] , SWIT_wire, \SADR/pgaddwy[17] , 
        \SADR/pgaddxz[2] , \REGF/RI_TBAI[10] , \REGF/RO_SRDA[7] , \pk_pc_h[1] , 
        \CODEIF/n3999 , \CODEQ/nqueue1[1] , \ALUIS/n3744 , \PDOSEL/n99 , 
        \CODEQ/nqueue2[2] , \ph_segset_h[18] , \BLU/n1587 , \pk_pdo_h[2] , 
        \stream4[25] , \SADR/pgaddxy[1] , \pgldi[21] , \SADR/pgaddyz[8] , 
        \pk_indy_h[0] , \pk_s3ba_h[9] , \pk_saba_h[15] , \stream4[16] , 
        \stream4[0] , \REGF/RI_PCOL[7] , \pgldi[12] , \REGF/RO_LLPSAS[1] , 
        \LBUS/n1392 , \LBUS/n1413 , \pk_s6ba_h[5] , ph_lbe2_h, 
        \REGF/RO_SRDA[20] , \PDOSEL/n106 , \BLU/n1479 , \pk_idcz_h[6] , 
        \MAIN/b_exec_stage , \CODEQ/nqueue1[50] , \ADOSEL/n4133 , 
        \CODEIF/n4030 , \CODEQ/nqueue1[49] , \REGF/RO_SRDA[13] , 
        \REGF/RO_PPCN[16] , \REGF/n8175 , \pkdptout[6] , \REGF/pk_indw_h[28] , 
        \REGF/n8152 , pkaccovf, pk_excp_h, \pk_s8ba_h[0] , \pk_sbba_h[14] , 
        \REGF/pk_indw_h[31] , \poalufnc[0] , \CODEIF/pgfpcel169 , 
        \CODEQ/nqueue2[39] , \CODEQ/nqueue2[20] , \ALUSHT/pkaluout[20] , 
        \CODEIF/pfctr[0] , \CODEIF/n3867 , \LBUS/n1434 , \CODEQ/nqueue2[13] , 
        \PDOSEL/n121 , \CODEIF/n4017 , \pgld16[8] , \ALUSHT/pkaluout[13] , 
        \SADR/pgaddwyz[20] , \pk_s4ba_h[12] , \pk_saba_h[8] , \ph_segset_h[9] , 
        \pk_saco_lh[21] , \ADOSEL/n4114 , \pk_sati_h[2] , \CODEIF/pfctr[16] , 
        \pk_sdba_h[4] , \LDIS/n3128 , \CONS/n600 , \BLU/n1562 , pktblcendh, 
        \REGF/RO_PCON[6] , \pk_saco_lh[12] , \pk_dpr_h[6] , 
        \SADR/pgaddwyz[13] , \pk_ada_h[3] , \CONS/n530 , \SADR/pgaddwxyz[2] , 
        \pk_indx_h[16] , \MAIN/n3625 , pk_sasea_h, \REGF/RI_SPR[24] , 
        \LBUS/ilt[2] , \ph_cpudout[29] , \ph_cpudout[30] , \SADR/lmtaddr[5] , 
        \pgldi[0] , \pk_rwrit_h[11] , \REGF/RI_SPR[17] , \pk_rwrit_h[22] , 
        \CODEIF/pgctrinc[3] , \pkbludgh[12] , \BLU/n1545 , \pk_rread_h[42] , 
        \CONS/n627 , \SADR/pgaddxy[17] , \SADR/pgaddwxyz[14] , \pk_pdo_h[18] , 
        \stream1[0] , \CONS/n612 , \pk_pcs2_h[12] , \pk_idcz_h[17] , 
        \CODEIF/n3949 , \BLU/n1570 , \pk_spr_h[23] , \pk_spr_h[10] , 
        \pk_sra1_h[21] , \pk_sra1_h[12] , \pk_sra2_h[0] , \SADR/pgaddwxz[22] , 
        \SADR/pgaddwxz[11] , \pk_s3ba_h[13] , \REGF/RI_TBAI[2] , 
        \REGF/RO_PPCN[6] , \ph_pdis_h[8] , \SAEXE/sequen , \CONS/n522 , 
        \LDCHK/n3234 , \LBUS/nlt[4] , \REGF/RO_EST1[2] , \ph_segset_h[26] , 
        \REGF/RO_EST2[1] , \MAIN/sprw_inhibith , \MAIN/n3610 , 
        \ALUSHT/pkshtout[23] , \MAIN/ph_rdwr2selh , \ph_segset_h[15] , 
        \pk_rwrit_h[0] , \pk_pcs2_h[0] , \stream4[31] , \CONS/n635 , 
        \stream4[28] , \ALUSHT/pkshtout[10] , \CODEIF/n3852 , \LDCHK/lpex[1] , 
        \PDOSEL/n114 , \BLU/n1557 , \LBUS/n1591 , \CONS/n699 , \CONS/n709 , 
        \SADR/pgaddwz[1] , \pk_indx_h[2] , \pk_s2ba_h[3] , \REGF/RO_ERRA[5] , 
        \CODEIF/n4022 , \LBUS/n1401 , \pgmuxout[6] , \ADOSEL/n4121 , 
        \REGF/RI_ACC[7] , \REGF/n8167 , \MAIN/ovferlth , \PDOSEL/n224 , 
        \pk_seba_h[15] , \REGF/RI_SRDA[11] , \REGF/RI_ACC[30] , 
        \REGF/RI_ACC[29] , \LDCHK/n3298 , \LDCHK/n3308 , \REGF/n8140 , 
        \SAEXE/srcrd_st , \SADR/pgaddwy[2] , \SADR/m_fadrl[17] , 
        \pgregadrh[1] , \CODEIF/n3875 , \LBUS/n1426 , \PDOSEL/n133 , 
        \REGF/RI_SRDA[22] , \ADOSEL/n4096 , \LDIS/ldexch[26] , \ADOSEL/n4106 , 
        \CODEIF/n4005 , \ALUIS/n3738 , \SADR/pgaddwxyz[19] , \SADR/lmtaddr[8] , 
        \pk_saba_h[5] , \pk_sdba_h[9] , \REGF/RI_PCOH[20] , 
        \REGF/RI_SRA12M[7] , \stream3[43] , wexacc, \pk_ada_h[13] , 
        \stream1[20] , \CONS/SACO[1] , \ph_cpudout[6] , \pk_sfba_h[14] , 
        \LBUS/n1448 , \CONS/n740 , \pk_ada_h[20] , \REGF/RI_EACC[6] , 
        \REGF/RI_PCOH[13] , \pgld32[3] , \stream1[13] , \pk_rread_h[56] , 
        \REG_2/n436 , \pk_pdo_h[15] , \pk_rwrit_h[36] , \pk_trba_h[23] , 
        \REGF/n8239 , \ph_cpudout[17] , \pk_spr_h[19] , \pk_dpr_h[2] , 
        \pk_trba_h[19] , \pk_trba_h[10] , \pk_pdo_h[26] , \REGF/n8099 , 
        \REGF/n8109 , \SADR/pgaddwx[23] , \SADR/pgaddwx[10] , 
        \SADR/pgaddyz[5] , \SADR/pgaddxyz[17] , \pk_indw_h[21] , 
        \pk_stat_h[1] , stage_2, \REG_2/RETCNT[6] , \ph_cpudout[24] , 
        \pgaluinb[21] , ph_word16h, \pk_indw_h[12] , \pk_s3ba_h[4] , 
        \pk_s6ba_h[8] , polcore_end, \pgaluinb[12] , \CODEQ/nqueue1[44] , 
        ph_byrtendh, \CODEIF/n3890 , \CODEIF/n3900 , \pgld16[5] , \BLU/n1539 , 
        \ph_segset_h[4] , \REGF/RI_PCOL[22] , \CODEIF/n3927 , \LDIS/n3154 , 
        \pk_indy_h[16] , \pk_s0ba_h[12] , \REGF/RI_PCOL[11] , 
        \REGF/RI_EACC[11] , \REGF/RI_EACC[22] , \CODEQ/nqueue2[34] , 
        \SADR/pgaddwxyz[23] , \SADR/pgaddwxyz[6] , \pk_s9ba_h[14] , 
        \REGF/n8182 , \REG_2/ph_retcnt_h[4] , \pk_rwrit_h[15] , 
        \REGF/pk_indw_h[25] , \REGF/n8199 , \pgldi[4] , \CONS/n346 , 
        \CONS/n557 , \SAEXE/n427 , \SADR/pgaddwxyz[10] , \pk_indx_h[12] , 
        \REGF/RI_SPR[20] , \LDCHK/n3266 , rmw22, \CONS/n667 , 
        \SADR/lmtaddr[1] , \pk_rread_h[46] , ph_tprsel_h, \SADR/pgaddwyz[17] , 
        \pk_indx_h[21] , \REGF/RI_SPR[13] , \pk_rwrit_h[26] , \BLU/n1505 , 
        \CODEIF/pgctrinc[7] , \BLU/n1495 , \pk_s4ba_h[16] , \pk_ada_h[30] , 
        \pk_ada_h[29] , \ALUIS/n3671 , \CONS/n640 , \BLU/n1522 , 
        \REGF/pk_indx_h[25] , \CODEIF/pfctr[12] , \SAEXE/stage_2nd , 
        \pk_sdba_h[0] , \pk_saco_lh[16] , \pk_ada_h[7] , \CONS/SACO[8] , 
        \CONS/n570 , \LDCHK/n3241 , \REGF/RO_PCON[2] , \REGF/RI_PCOL[18] , 
        \poalufnc[4] , \CODEIF/pfctr[4] , \SADR/pgaddwx[19] , \pk_indy_h[4] , 
        \poshtfnc[1] , \ALUSHT/pkaluout[24] , \CODEIF/n3765 , 
        \CODEQ/nqueue2[24] , \pk_s8ba_h[4] , \REGF/n8082 , \REGF/n8112 , 
        \ADOSEL/n4154 , \ALUSHT/pkaluout[17] , \pk_sbba_h[10] , 
        \REGF/RI_EACC[18] , \REGF/n8222 , \CODEQ/nqueue2[17] , \PDOSEL/n161 , 
        \SADR/pgaddwy[20] , \SADR/pgaddwy[13] , \SADR/pgaddxy[5] , 
        \pk_s6ba_h[1] , ph_tcer_h, \REGF/RO_SRDA[24] , \pk_idcz_h[2] , 
        \REGF/n8205 , \CODEIF/n3990 , \CODEQ/nqueue1[54] , \PDOSEL/n146 , 
        \REGF/RO_SRDA[17] , \REGF/RO_PSASH[15] , \REGF/RO_LLPSAS[5] , 
        \LBUS/n1453 , \REGF/RO_PPCN[12] , \pgaluinb[28] , \pgaluinb[31] , 
        \MAIN/st_swctl , \REGF/pk_indy_h[31] , \REGF/pk_indy_h[28] , 
        \pkdptout[2] , \LBUS/access_en_h , \REGF/n8135 , ph_lwdsrch, 
        \pgldi[25] , \MAIN/EXCEP_1H , \SADR/pgaddxz[6] , \pk_rwrit_h[9] , 
        \MAIN/a_exec_stage , \REGF/pk_idcz_h[29] , \ALUIS/n3723 , 
        \pk_pcs2_h[9] , phlbdir, \REGF/pk_idcz_h[30] , \pk_pdo_h[6] , 
        \stream4[38] , \stream4[21] , \ALUSHT/pkshtout[19] , \CONS/n735 , 
        ph_cperr_h, \PDOSEL/n128 , \CMPX/n1050 , \SADR/pgaddwxz[18] , 
        \pk_saba_h[11] , \REGF/RI_PCOL[3] , \stream4[12] , \pgldi[16] , 
        \CONS/n595 , \stream4[4] , \LDCHK/n3283 , \LDCHK/n3313 , \RSTGN/n_6 , 
        \pgsdprhh[31] , \pgsdprhh[28] , \ph_pdis_h[1] , \pk_sra1_h[31] , 
        \pk_sra1_h[28] , \SADR/pgovfwyz , \pk_seba_h[7] , \REGF/RO_SRDA[3] , 
        oltff, \SAEXE/adovflth1 , \stream1[9] , \CODEQ/nqueue2[6] , 
        \pk_pc_h[5] , \CODEIF/n4039 , \ALUIS/n3694 , \ALUIS/n3704 , 
        \UPIF/iready , \CODEQ/nqueue1[5] , \CONS/n682 , \CONS/n712 , 
        \REGF/RI_TBAI[14] , \CODEIF/n3849 , \BLU/n1470 , \pgregadrh[8] , 
        \pk_s9ba_h[3] , \CODEIF/n3975 , \PDOSEL/n75 , \pk_pc_h[13] , 
        \REGF/RI_DPR[21] , \stream3[53] , \pgld16[11] , \SADR/pgaddwz[8] , 
        \REGF/RI_SRDA[18] , \REGF/RO_LPSAS2156[11] , \pk_indw_h[6] , 
        \pk_s7ba_h[17] , \REGF/pk_seba_h[18] , \REGF/RI_DPR[12] , 
        \LDCHK/pglpinff[1] , \pk_s7ba_h[6] , \REGF/RO_EACC[24] , \CONS/n539 , 
        \REGF/pk_stat_h[31] , \REGF/RI_STAT[1] , \REGF/n8067 , \pk_sra2_h[9] , 
        \SADR/segbase[4] , \REGF/RO_EACC[17] , \REGF/RI_ACC[20] , 
        \CODEIF/n3952 , phrelbsth, \CONS/n609 , \SADR/pgaddxy[16] , 
        \SADR/pgaddwxz[23] , \SADR/pgaddwxz[10] , \pk_s3ba_h[12] , 
        \ph_segset_h[27] , \REGF/RO_EST2[0] , \LDIS/n3121 , \REGF/RI_ACC[13] , 
        \ALUSHT/pkshtout[22] , \ph_segset_h[14] , \REGF/RI_TBAI[3] , 
        \REGF/RO_EST1[3] , \stream4[30] , \stream4[29] , \ALUSHT/pkshtout[11] , 
        \CONS/n625 , \BLU/n1547 , \pk_rwrit_h[1] , \pk_pcs2_h[1] , 
        \CODEIF/n3959 , \CONS/n602 , \BLU/n1560 , \REGF/RO_PPCN[7] , 
        \stream1[1] , \stream2[2] , \BLU/SRC_DATA_M , \ph_pdis_h[9] , 
        pgldperrh, \MAIN/n3627 , \LBUS/nlt[5] , \pk_idcz_h[16] , \CONS/n532 , 
        n10737, \pk_spr_h[22] , \pk_spr_h[11] , \pk_sra1_h[20] , 
        \pk_sra1_h[13] , ph_cperlt_h, \pk_pcs2_h[13] , \SAEXE/seq_end , 
        \SADR/pgaddwy[3] , \SADR/pgaddwz[0] , \REGF/RI_SRDA[10] , \REGF/n8150 , 
        \stream3[42] , \ADOSEL/n4116 , \CODEIF/n4015 , \ALUIS/n3728 , 
        \pk_sra2_h[1] , \SADR/m_fadrl[16] , \CODEIF/n3865 , ph_bnolt_h, 
        \PDOSEL/n123 , \LDIS/ldexch[27] , \pk_s2ba_h[2] , \pgregadrh[0] , 
        \REGF/RI_SRDA[23] , \LBUS/n1436 , \REGF/RO_ERRA[4] , \pgmuxout[7] , 
        \REGF/RI_ACC[6] , \ADOSEL/n4131 , \CODEIF/n4032 , \CODEIF/n3842 , 
        \LDCHK/lpex[0] , \LBUS/n1411 , \PDOSEL/n104 , \CONS/n719 , 
        \pk_trba_h[22] , \pk_indx_h[3] , \pk_seba_h[14] , ph_ovfihbh, 
        \CONS/n689 , \REGF/RI_ACC[28] , \LDCHK/n3288 , \REGF/RI_ACC[31] , 
        \REGF/n8177 , \ph_cpudout[16] , \SADR/pgaddwxyz[18] , 
        \SADR/lmtaddr[9] , \pk_rread_h[57] , \pk_pdo_h[14] , \REGF/n8229 , 
        \pk_trba_h[11] , \pk_rwrit_h[37] , \ph_cpudout[25] , \BLU/n1585 , 
        \REGF/n8089 , \REGF/n8119 , ph_ioselh, \REG_2/RETCNT[7] , 
        \pk_dpr_h[3] , \pk_trba_h[18] , \SADR/pgaddwx[22] , \SADR/pgaddwx[11] , 
        \SADR/pgovfxyz , \pk_sdba_h[8] , \REGF/RI_PCOH[21] , \pk_pdo_h[27] , 
        obacc, \stream1[21] , \ph_cpudout[7] , \pk_ada_h[12] , 
        \LBUS/ph_lbusylth , \pk_indy_h[17] , \pk_s0ba_h[13] , \pk_saba_h[4] , 
        \REGF/RI_SRA12M[6] , \REGF/RI_EACC[7] , \pgld32[2] , \CONS/SACO[0] , 
        \pk_sfba_h[15] , \REGF/RI_PCOH[12] , \stream1[12] , \ALUIS/n3746 , 
        \pk_ada_h[21] , seg_cnfg_h, \LBUS/n1458 , \REGF/RI_EACC[10] , 
        \CODEIF/n3937 , \SADR/pgaddyz[4] , \LDIS/n3144 , \SADR/pgaddxyz[16] , 
        \ph_segset_h[5] , \REGF/RI_PCOL[23] , \pgld16[4] , \SADR/pgaddwyz[16] , 
        \pk_indw_h[20] , \pk_s9ba_h[15] , \REGF/pk_indw_h[24] , 
        \REGF/RI_EACC[23] , \CODEQ/nqueue2[35] , \REGF/RI_PCOL[10] , phsaerrh, 
        \REGF/n8192 , \REG_2/ph_retcnt_h[5] , cf_wait, cnfg_write_h, 
        \pk_indw_h[13] , \pk_s6ba_h[9] , \pk_stat_h[0] , \pgaluinb[20] , 
        \BLU/n1529 , \pk_s3ba_h[5] , \CODEIF/n3880 , \pk_s4ba_h[17] , 
        \CODEIF/pfctr[13] , \CODEIF/n3910 , \pgaluinb[13] , \LDIS/n3163 , 
        \MAIN/LBAOVFH , \CODEQ/nqueue1[45] , \pk_sdba_h[1] , \pk_saco_lh[17] , 
        \REGF/pk_indx_h[24] , \pk_ada_h[31] , \CONS/n650 , \pk_ada_h[28] , 
        \BLU/n1532 , \LDCHK/n3251 , \REGF/RO_PCON[3] , \SADR/pgovfwx , 
        \pk_indx_h[13] , \pk_ada_h[6] , \CONS/SACO[9] , \CONS/n560 , 
        \REGF/RI_SPR[21] , \LDCHK/n3276 , \SADR/pgaddwxyz[22] , 
        \pk_rwrit_h[14] , \REGF/n8189 , ph_piosl_h, \CONS/n547 , 
        \SADR/pgaddwxyz[7] , \pgldi[5] , \pk_indx_h[20] , \CODEIF/pgctrinc[6] , 
        \ALUIS/n3661 , \SADR/lmtaddr[0] , \REGF/RI_SPR[12] , \pk_rread_h[47] , 
        \REGF/pk_sfba_h[18] , \CONS/n677 , \SADR/pgaddwxyz[11] , 
        \pk_rwrit_h[27] , \BLU/n1485 , \pgsdprhh[30] , \pgsdprhh[29] , 
        \pk_spr_h[18] , \BLU/n1515 , \SADR/pgaddwx[18] , \pk_indy_h[5] , 
        \pk_s6ba_h[0] , \REGF/RO_SRDA[25] , \REGF/n8215 , \CODEIF/n3980 , 
        \pk_idcz_h[3] , \REGF/RO_LLPSAS[4] , \LBUS/n1443 , \PDOSEL/n156 , 
        \PDOSEL/n80 , \CODEQ/nqueue1[55] , \REGF/pk_indy_h[30] , 
        \REGF/pk_indy_h[29] , \pkdptout[3] , \REGF/pk_s9ba_h[18] , 
        \REGF/RO_SRDA[16] , \REGF/RO_PPCN[13] , \REGF/n8125 , \REGF/n8102 , 
        \poshtfnc[0] , \pgaluinb[29] , ph_srdalth, \pgaluinb[30] , 
        \CODEQ/nqueue2[25] , \REGF/n8092 , \REGF/RI_PCOL[19] , \REGF/n8232 , 
        \CODEIF/pfctr[5] , \ALUSHT/pkaluout[25] , phlmterrh, \pk_s8ba_h[5] , 
        \pk_sbba_h[11] , \REGF/RI_EACC[19] , \ADOSEL/n4144 , 
        \ALUSHT/pkaluout[16] , \CODEQ/nqueue2[16] , \pk_seba_h[6] , 
        \ph_pdis_h[0] , \LDCHK/n3293 , \LDCHK/n3303 , pgrstith, \pk_spr_h[15] , 
        \pk_sra1_h[30] , \pk_sra2_h[8] , \SADR/pgaddwy[21] , 
        \SADR/pgaddwy[12] , \SADR/pgaddxz[7] , \SADR/pgovfwxz , 
        \REGF/RI_TBAI[15] , \pk_pc_h[4] , \CONS/n702 , \CODEQ/nqueue1[4] , 
        \CONS/n692 , \REGF/RO_SRDA[2] , \CODEIF/n3859 , \CODEIF/n4029 , 
        \ALUIS/n3684 , \ALUIS/n3714 , \CODEQ/nqueue2[7] , \pk_pdo_h[7] , 
        \stream4[20] , \ALUSHT/pkshtout[18] , \CONS/n725 , \stream4[39] , 
        \PDOSEL/n138 , po_brsel_h, \SADR/pgaddxy[4] , \pgldi[24] , 
        \SADR/pgaddwxz[19] , \pk_saba_h[10] , \pk_rwrit_h[8] , \pk_pcs2_h[8] , 
        \REGF/pk_idcz_h[31] , \REGF/pk_idcz_h[28] , ph_aluovf_h, \ALUIS/n3733 , 
        \stream4[13] , \REGF/RI_PCOL[2] , \stream4[5] , \CONS/n585 , 
        \pgldi[17] , \SADR/segbase[5] , \pk_s7ba_h[7] , \REGF/pk_stat_h[30] , 
        \REGF/RI_ACC[21] , \pk_s7ba_h[16] , \CONS/n338 , \REGF/RO_EACC[25] , 
        \REGF/RI_STAT[0] , \REGF/n8077 , \CONS/n529 , \MAIN/single_write , 
        \REGF/RI_ACC[12] , \REGF/RO_EACC[16] , ciffsel, \CODEIF/n3942 , 
        \LDIS/n3131 , \pk_pc_h[12] , \REGF/RI_DPR[20] , \CONS/n619 , 
        \pk_sra1_h[29] , \SADR/pgaddwx[15] , \SADR/pgaddwz[9] , \pgregadrh[9] , 
        \pk_s9ba_h[2] , \stream3[52] , \CODEIF/n3965 , \pgld16[10] , 
        \REGF/RI_DPR[13] , \LDCHK/pglpinff[0] , \LDIS/n3116 , \SAEXE/srcread , 
        \SADR/pgaddyz[0] , \pk_indw_h[17] , \pk_indw_h[7] , \REGF/RI_SRDA[19] , 
        \REGF/RO_LPSAS2156[10] , \LBUS/n1606 , \pk_s3ba_h[1] , ph_sdirlth, 
        \REGF/pk_indy_h[24] , \REGF/n8065 , \CODEIF/fm_config[0] , 
        \pgaluinb[24] , \phshtd[2] , \REGF/RO_SRDA[31] , \REGF/RO_SRDA[28] , 
        \REGF/RO_LLPSAS[9] , \REGF/pk_sbba_h[18] , \pgaluinb[17] , 
        \CODEQ/nqueue1[41] , \CODEQ/nqueue1[58] , \CODEIF/n3950 , \LDIS/n3123 , 
        \BLU/n1569 , \pk_s8ba_h[8] , \REGF/RI_PCOL[27] , \REG_2/ncnt3[0] , 
        \pgld16[0] , \SADR/pgaddxyz[12] , \ph_segset_h[1] , 
        \SADR/pgaddxyz[21] , \pk_indy_h[13] , \pk_s0ba_h[17] , 
        \REGF/RI_EACC[14] , \CODEIF/n3977 , \PDOSEL/n77 , \pk_indy_h[20] , 
        \pk_indy_h[8] , \pk_s9ba_h[11] , \REGF/RI_PCOL[14] , 
        \ALUSHT/pkaluout[31] , \ALUSHT/pkaluout[28] , \CODEIF/pfctr[8] , 
        stage_a, \REG_2/ph_retcnt_h[1] , \pk_saba_h[0] , \pk_sfba_h[11] , 
        \REGF/RI_PCOH[25] , \REGF/RI_SRA12M[2] , \REGF/RI_EACC[27] , ph_sais_h, 
        \CODEQ/nqueue2[28] , \UPIF/alusfterr , \CODEQ/nqueue2[31] , 
        \CONS/SACO[4] , \pk_ada_h[16] , \stream1[25] , \LDCHK/n3281 , 
        \LDCHK/n3311 , \ph_cpudout[3] , \pk_ada_h[25] , \LBUS/n1399 , 
        \LBUS/n1418 , \CONS/n680 , \BLU/n1472 , \CONS/n710 , 
        \REGF/RI_PCOH[16] , \REGF/pk_indx_h[30] , \REGF/pk_indx_h[29] , 
        \ADOSEL/n4138 , \REGF/RI_EACC[3] , \ALUIS/n3696 , \ALUIS/n3706 , 
        \pk_rwrit_h[33] , \pgld32[6] , \pgldi[8] , ph_tblcdech, 
        \pk_rread_h[53] , \REGF/n8269 , \pk_pdo_h[10] , \ALUIS/n3721 , 
        \CONS/n737 , \ph_cpudout[12] , \pk_rread_h[60] , \pk_pdo_h[23] , 
        \CONS/n597 , \pk_rwrit_h[19] , \REGF/n8159 , \REG_2/RETCNT[3] , 
        \pk_sra1_h[17] , \pk_sra2_h[5] , \pk_trba_h[15] , \LBUS/n1451 , 
        \ph_cpudout[21] , \PDOSEL/n92 , \SADR/pgaddwy[7] , \SADR/pgaddwz[4] , 
        \pk_indx_h[7] , \SADR/segbase[8] , \pk_s2ba_h[6] , \REGF/n8207 , 
        \PDOSEL/n144 , \CODEIF/n3992 , ph_adrinc_h, \REGF/RO_ERRA[0] , 
        \REGF/RI_ACC[2] , \pgmuxout[3] , \REGF/RO_EACC[31] , \REGF/n8137 , 
        \REGF/RO_EACC[28] , \LBUS/temp[3] , \pk_seba_h[10] , \REGF/n8080 , 
        po_sprlth, \REGF/n8110 , \SADR/m_fadrl[21] , \REGF/RI_SRDA[14] , 
        \SADR/m_fadrl[12] , \pgregadrh[4] , \SADR/intbitno[1] , 
        \REGF/RI_SRDA[27] , \REGF/n8220 , \LDIS/ldexch[23] , pgoddflgh, 
        \stream3[46] , \PDOSEL/n163 , pktrscovfh, \ADOSEL/n4156 , 
        \pk_idcz_h[21] , \SADR/pgaddxy[12] , \REGF/RI_TBAI[18] , \BLU/n1520 , 
        \pk_pc_h[9] , \CODEIF/n3889 , \CODEIF/n3919 , \LDIS/ldexcl[12] , 
        pgbnolth, \CONS/n642 , \pk_pcs2_h[17] , \CODEQ/nqueue1[9] , step2_cf, 
        \SADR/pgaddwy[16] , \SADR/pgaddxy[21] , \REGF/RO_PPCN[3] , 
        \pk_idcz_h[12] , \LDCHK/n3243 , \CONS/n572 , 
        \LBUS/*cell*3982/U111/CONTROL2 , \LBUS/*cell*3982/U176/CONTROL1 , 
        \LBUS/nlt[1] , \SADR/pgaddxy[9] , \SADR/pgaddwxz[14] , \pk_s3ba_h[16] , 
        \REGF/RI_TBAI[7] , \REGF/RO_EST1[7] , \pgbitnoh[2] , \ph_segset_h[23] , 
        \stream4[8] , po_bitsrc_h, \SAEXE/n425 , \LDCHK/n3264 , 
        \ALUSHT/pkshtout[26] , \CONS/n344 , \pk_rwrit_h[5] , \pk_pcs2_h[5] , 
        \REGF/pk_idcz_h[25] , \CONS/n555 , \pgldi[30] , \ALUIS/n3673 , 
        \SADR/pgaddxy[0] , \pk_indw_h[3] , \pk_s9ba_h[6] , \ph_segset_h[10] , 
        \pgldi[29] , \BLU/n1497 , \BLU/n1507 , \stream4[34] , \CONS/n665 , 
        \LDIS/n3156 , \ALUSHT/pkshtout[15] , \pk_pc_h[16] , \stream3[56] , 
        \CODEIF/n3925 , \pgld16[14] , \ALUIS/n3668 , \REGF/RI_DPR[24] , 
        \REGF/n8180 , \SADR/segbase[1] , \pk_s7ba_h[12] , \REGF/RO_EACC[21] , 
        \REGF/RI_DPR[17] , \LDIS/ldexch[19] , phbnolth, \REGF/RI_STAT[4] , 
        \SAEXE/wrd_datah , \LDCHK/n3258 , \CONS/n569 , \SAEXE/n419 , 
        \pk_s7ba_h[3] , \REGF/RI_ACC[25] , \REGF/RO_ERRA[9] , 
        \REGF/RO_EACC[12] , \CODEIF/n3892 , \CODEIF/n3902 , \CONS/n659 , 
        \REGF/RI_ACC[16] , \pgldi[20] , \SADR/pgaddxz[3] , \pk_saba_h[14] , 
        \ph_segset_h[19] , \pk_pdo_h[3] , \PDOSEL/n178 , \stream4[24] , 
        \REGF/RI_PCOL[6] , \pgldi[13] , \stream4[17] , \stream4[1] , phrstihb, 
        phrstith, \SADR/pgaddyz[9] , \pk_indy_h[1] , \pk_seba_h[2] , 
        \REGF/RI_TBAI[22] , \ph_pdis_h[4] , \REGF/RI_TBAI[11] , 
        \REGF/RO_SRDA[6] , \CODEQ/nqueue2[3] , \CODEIF/n3989 , \ALUIS/n3754 , 
        \pk_pc_h[0] , \REGF/pk_indw_h[30] , \poalufnc[1] , \CODEIF/pfctr[1] , 
        \ALUSHT/pkaluout[21] , \CODEQ/nqueue1[0] , \CONS/n742 , \CMPX/n1049 , 
        \REGF/pk_indw_h[29] , \pk_s8ba_h[1] , \REGF/n8142 , 
        \CODEQ/nqueue2[38] , \CODEQ/nqueue2[21] , \pk_sbba_h[15] , 
        \ADOSEL/n4094 , \ph_segset_h[8] , \pk_idcz_h[7] , \ADOSEL/n4104 , 
        \CODEIF/n3877 , \CODEIF/n4007 , \ALUSHT/pkaluout[12] , \pgld16[9] , 
        \LBUS/n1424 , \CODEQ/nqueue2[12] , \CODEIF/n4020 , \PDOSEL/n131 , 
        \REGF/RO_LLPSAS[0] , \ADOSEL/n4123 , \CODEQ/nqueue1[51] , 
        \CODEQ/nqueue1[48] , \LBUS/n1403 , \LBUS/n1593 , \PDOSEL/n116 , 
        \BLU/n1469 , \pk_dpr_h[7] , \SADR/pgaddwxyz[15] , \SADR/pgaddwxyz[3] , 
        \pk_s3ba_h[8] , \REGF/RO_SRDA[21] , \CODEIF/n3850 , \pk_s6ba_h[4] , 
        \REGF/RO_SRDA[12] , \REGF/RO_PPCN[17] , \REGF/n8165 , \PDOSEL/n226 , 
        \pgldi[1] , \pkdptout[7] , \pk_indx_h[17] , \pk_rwrit_h[10] , 
        ph_dprsel2_h, \REGF/RI_SPR[25] , \REGF/n8059 , \MAIN/n3612 , 
        \LDCHK/n3236 , \ph_cpudout[28] , \ph_cpudout[31] , \pk_rwrit_h[23] , 
        \BLU/n1555 , \pk_pdo_h[19] , \CONS/n637 , \pk_dpr_h[5] , 
        \SADR/pgaddwyz[21] , \SADR/lmtaddr[4] , \pk_rread_h[43] , 
        \REGF/RI_SPR[16] , \CODEIF/pgctrinc[2] , \pkbludgh[13] , \BLU/n1572 , 
        \SADR/pgaddwyz[12] , \pk_s4ba_h[13] , \pk_saco_lh[20] , \LDIS/n3138 , 
        \CONS/n610 , \CODEIF/pfctr[17] , pkshterr, \pk_saba_h[9] , 
        \pk_ada_h[2] , \CONS/n520 , \SADR/pgaddxyz[19] , \pk_indy_h[18] , 
        \pk_indy_h[3] , \pk_sdba_h[5] , \REGF/RO_PCON[7] , \pk_saco_lh[13] , 
        \REGF/n8162 , \CODEQ/nqueue2[23] , srctype0, \poalufnc[3] , 
        \CODEIF/pfctr[3] , \MAIN/dprw_tap2 , \CODEIF/n3857 , 
        \ALUSHT/pkaluout[23] , \PDOSEL/n111 , \ADOSEL/n4124 , \CODEIF/n4027 , 
        \LBUS/n1404 , \CODEQ/nqueue2[10] , \LBUS/n1594 , \ALUSHT/pkaluout[10] , 
        \SADR/pgaddwxyz[17] , \SADR/pgaddwxyz[1] , \pk_indx_h[15] , 
        \pk_s6ba_h[6] , \pk_s8ba_h[3] , \pk_sbba_h[17] , \REGF/RO_SRDA[23] , 
        \pk_idcz_h[5] , \REGF/pk_s0ba_h[18] , \CODEIF/n3870 , ph_word32h, 
        \PDOSEL/n136 , \ADOSEL/n4103 , \LBUS/n1423 , \pkdptout[5] , 
        \ADOSEL/n4093 , \CODEQ/nqueue1[53] , \CODEIF/n4000 , ph_lbe1_h, 
        \REGF/RO_SRDA[10] , \REGF/n8145 , \REGF/RO_PPCN[15] , 
        \REGF/RI_SPR[27] , \pgldi[3] , \pk_rwrit_h[12] , \REGF/n8079 , 
        \LBUS/ilt[1] , \MAIN/n3632 , \pk_pdo_h[31] , \pk_pdo_h[28] , 
        \CONS/n527 , \SADR/lmtaddr[6] , \REGF/RI_SPR[14] , 
        \CODEIF/pgctrinc[0] , \pkbludgh[11] , \ph_cpudout[19] , 
        \pk_rread_h[41] , po_raccen_h, \pk_rread_h[58] , \pk_s4ba_h[11] , 
        \pk_rwrit_h[38] , \CONS/n617 , \BLU/n1575 , \pk_rwrit_h[21] , 
        \CODEIF/pfctr[15] , \REGF/RO_EST2[15] , \REGF/RI_EACC[8] , 
        \SAEXE/sa_start3 , \pk_saco_lh[22] , \LDIS/n3118 , \CONS/n630 , 
        ph_oprtrs_h, \SADR/pgaddwyz[23] , \pk_sati_h[1] , \SADR/pgaddwyz[10] , 
        \pk_sdba_h[7] , \pk_saco_lh[11] , ph_lbaovf, \BLU/n1552 , 
        \LDCHK/n3231 , \ph_cpudout[8] , \REGF/RO_PCON[5] , \REGF/RI_SRA12M[9] , 
        ph_timsth, \pk_indw_h[1] , \SADR/m_fadrl[19] , \pk_s9ba_h[4] , 
        \pk_pc_h[14] , \pk_ada_h[0] , \MAIN/n3615 , \REGF/RI_DPR[26] , 
        \LBUS/n1608 , \pk_stat_h[18] , \stream3[54] , \CODEIF/n3895 , 
        \CODEIF/n3905 , \LDIS/ldexch[31] , \REGF/RI_DPR[15] , 
        \LDIS/ldexch[28] , \SADR/segbase[3] , \pk_s7ba_h[1] , 
        \REGF/RI_ACC[27] , ph_extselh, \LDCHK/n3278 , \pk_s7ba_h[10] , 
        \CONS/n549 , \REGF/RO_EACC[23] , \REGF/n8187 , \REGF/RO_EACC[10] , 
        \REGF/RI_ACC[14] , \pgmuxout[8] , \REGF/RI_ACC[9] , \pk_pdo_h[1] , 
        \CODEIF/n3922 , \LDIS/n3151 , \CONS/n679 , \CONS/n745 , 
        \SADR/pgaddwy[14] , \SADR/pgaddxz[1] , \stream4[26] , \PDOSEL/n158 , 
        \SADR/pgaddxy[2] , \pk_saba_h[16] , \pgldi[22] , \ALUIS/n3753 , 
        st_exectl, \LBUS/lnsa_err , \pk_seba_h[0] , \ph_segset_h[31] , 
        \ph_segset_h[28] , \stream4[15] , \stream4[3] , \pgldi[11] , 
        \REGF/RI_PCOL[4] , \MAIN/astregw_tap1 , \REGF/RI_TBAI[20] , 
        \ph_pdis_h[6] , \REGF/RO_PPCN[8] , \pk_idcz_h[19] , \SADR/m_fadrh[31] , 
        \SADR/m_fadrh[28] , \SADR/pgaddxy[19] , \pk_pc_h[2] , 
        \CODEQ/nqueue1[2] , \REGF/RI_TBAI[13] , \pk_sra1_h[15] , 
        \pk_sra2_h[7] , \pk_s2ba_h[4] , \REGF/RO_SRDA[4] , ph_ldaoutenhp, 
        \CODEQ/nqueue2[1] , \REGF/RO_ERRA[2] , \ADOSEL/n4151 , \pgmuxout[1] , 
        \REGF/RI_ACC[0] , \REGF/RO_EACC[19] , \REGF/n8227 , wonly2, 
        \PDOSEL/n164 , \pk_indx_h[5] , \pk_s7ba_h[8] , \pk_seba_h[12] , 
        \REGF/n8087 , \REGF/n8117 , \SADR/pgaddwy[5] , \REGF/pk_sctio_h , 
        \SADR/pgaddwz[6] , \SADR/m_fadrl[23] , \SADR/pgaddxy[10] , 
        \pk_indw_h[8] , \REGF/RI_SRDA[16] , \REGF/n8130 , \SADR/m_fadrl[10] , 
        \SADR/intbitno[3] , \stream3[44] , \ALUIS/n3748 , \REGF/RI_SRDA[25] , 
        \REGF/n8200 , \PDOSEL/n143 , \CODEIF/n3995 , \pgregadrh[6] , 
        \LDIS/ldexch[21] , \LBUS/n1456 , \PDOSEL/n95 , \CODEIF/n3939 , 
        \CONS/n662 , \LDIS/ldexcl[10] , phadrdech, \BLU/n1490 , \BLU/n1500 , 
        \CODEIF/friend_in , ph_dprtrs_h, \pk_idcz_h[23] , \CODEQ/nqueue2[8] , 
        \SADR/pgaddxy[23] , \ALUIS/n3674 , \pk_seba_h[9] , \REGF/RO_PPCN[1] , 
        \LBUS/nlt[3] , \CONS/n343 , \CONS/n552 , \pk_idcz_h[10] , 
        \LDCHK/n3263 , \SAEXE/n422 , \RSTGN/WRST_2H , \SADR/pgaddxz[8] , 
        \SADR/pgaddwxz[16] , \pgbitnoh[0] , \ph_segset_h[21] , 
        \REGF/RO_EST2[6] , \pk_pcs2_h[15] , \CONS/n575 , all0bsel, 
        \ALUSHT/pkshtout[24] , \LDCHK/n3244 , \pk_s3ba_h[14] , 
        \ph_segset_h[12] , \REGF/RI_TBAI[5] , \REGF/RO_EST1[5] , \pgldi[18] , 
        \pk_pdo_h[8] , \stream4[36] , \ALUSHT/pkshtout[17] , \CONS/n645 , 
        \BLU/n1527 , \REGF/RO_SRDA[19] , \pk_rwrit_h[7] , \ALUIS/n3653 , 
        \pk_pcs2_h[7] , \REGF/pk_idcz_h[27] , \REGF/pk_indy_h[26] , 
        \phshtd[0] , \pk_spr_h[17] , \SADR/pgaddwx[17] , \pk_indw_h[15] , 
        \pgaluinb[26] , \BLU/n1549 , \SAEXE/stage_1st , \pk_indy_h[11] , 
        \pk_s3ba_h[3] , \CODEIF/n3970 , \CODEIF/n3957 , \pgaluinb[15] , 
        \LBUS/*cell*3982/U70/CONTROL1 , \CODEQ/nqueue1[43] , \PDOSEL/n181 , 
        \pk_s0ba_h[15] , \REGF/RI_EACC[16] , \CODEQ/nqueue2[19] , \LDIS/n3124 , 
        \SADR/pgaddyz[2] , \ph_segset_h[3] , \SADR/pgaddwyz[19] , 
        \SADR/pgaddxyz[23] , \SADR/pgaddxyz[10] , \pk_indy_h[22] , 
        \REGF/RI_PCOL[25] , \pgld16[2] , \ALUSHT/pkaluout[19] , 
        \pk_s9ba_h[13] , \REGF/RI_EACC[25] , \CODEQ/nqueue2[33] , 
        \REG_2/ph_retcnt_h[3] , \REGF/RI_PCOL[16] , \REGF/n8062 , \MAIN/n3629 , 
        allfasel, \REGF/RI_PCOH[27] , \REGF/RI_SRA12M[0] , \pk_saco_lh[18] , 
        \stream1[27] , \pk_ada_h[14] , \ph_cpudout[1] , \pk_saba_h[2] , 
        \pk_ada_h[9] , \CONS/SACO[6] , \CONS/n590 , \pgld32[4] , 
        \pk_sfba_h[13] , \REGF/RI_PCOH[14] , \REGF/RI_EACC[1] , \stream1[14] , 
        \ALUIS/n3726 , \ADOSEL/n4088 , \ADOSEL/n4118 , \pk_ada_h[27] , 
        \LBUS/n1438 , \CONS/n730 , \CODEIF/pgctrinc[9] , \pk_rread_h[51] , 
        \pk_rread_h[48] , \pk_pdo_h[12] , \ALUIS/n3691 , \ALUIS/n3701 , 
        \ph_cpudout[10] , \CONS/n687 , \CONS/n717 , \pk_trba_h[17] , 
        \pk_rwrit_h[31] , \pk_rwrit_h[28] , \BLU/n1475 , \SADR/pgaddwxyz[8] , 
        \LDCHK/n3286 , \ph_cpudout[23] , \REGF/n8179 , \REG_2/RETCNT[1] , 
        \pk_rread_h[62] , \pk_pdo_h[21] , \pk_spr_h[30] , \pk_sra1_h[18] , 
        \SADR/pgaddwy[23] , \SADR/pgaddwy[10] , \SADR/pgaddxy[6] , 
        \SADR/pgovfyz , \pk_pcs2_h[18] , ph_tirtendh, \CMPX/n1047 , 
        \CONS/n582 , \SADR/sadr[0] , \pk_seba_h[4] , \ph_pdis_h[2] , 
        ph_sa1lt_h, \CODEIF/n3879 , \CODEIF/n4009 , \CODEQ/nqueue2[5] , 
        \ALUIS/n3734 , \REGF/RI_TBAI[17] , \pk_pc_h[6] , \stream2[9] , 
        \MAIN/ph_rrmwh , \ALUIS/n3683 , \ALUIS/n3713 , \CODEQ/nqueue1[6] , 
        \CONS/n722 , \pgldi[26] , \MAIN/EXCEP_2H , \SADR/pgaddxz[5] , 
        \PDOSEL/n118 , \BLU/n1467 , \pk_pdo_h[5] , \stream4[22] , ph_word32_h, 
        \CONS/n695 , \CONS/n705 , \SADR/pgaddwy[8] , \pk_indw_h[5] , 
        \pk_indx_h[8] , \SADR/segbase[7] , \pk_s7ba_h[14] , \pk_saba_h[12] , 
        \REGF/RI_PCOL[0] , \REGF/RI_TBAI[8] , \pgldi[15] , \LDCHK/n3294 , 
        \LDCHK/n3304 , \REGF/RO_EACC[27] , \stream4[11] , \stream4[7] , 
        \ALUSHT/pkshtout[29] , \ALUSHT/pkshtout[30] , \REGF/RI_STAT[2] , 
        \REGF/n8057 , \LBUS/n1601 , \REGF/RI_ACC[23] , \LDCHK/n3238 , 
        ph_bdstenh, \pk_s2ba_h[9] , \pk_s7ba_h[5] , \REGF/RO_EACC[14] , ronly1, 
        \CONS/n639 , \CODEIF/n3962 , \pk_s9ba_h[0] , \REGF/RI_SRDA[31] , 
        \REGF/RI_ACC[10] , \REGF/RI_SRDA[28] , \LDIS/n3136 , po_sprtrs_h, 
        \pk_pc_h[10] , \stream3[50] , \stream3[49] , \CODEIF/n3945 , 
        \pgld16[12] , \REGF/RI_DPR[22] , \REGF/n8070 , ph_lwdsrc_h, 
        \REGF/RI_DPR[11] , \SADR/pgaddwyz[14] , \pk_s4ba_h[15] , 
        \REGF/RI_PCOH[19] , \REGF/pk_indx_h[26] , \MAIN/cstregw_tap2 , 
        \LDCHK/pglpinff[2] , \LDIS/n3158 , \BLU/n1482 , \BLU/n1512 , 
        \CONS/n670 , \stream1[19] , \ALUIS/n3666 , \CODEIF/pfctr[11] , 
        \pgld32[9] , \pk_ada_h[19] , \pk_ada_h[4] , \CONS/n351 , \CONS/n540 , 
        ph_filewr_h, \SADR/pgaddwxyz[20] , \SADR/pgaddwxyz[5] , \pk_sdba_h[3] , 
        \pgldi[7] , \pk_saco_lh[15] , \REGF/RO_PCON[1] , \SAEXE/n430 , 
        \LDCHK/n3271 , \CONS/n567 , \pk_rwrit_h[16] , \pk_spr_h[29] , 
        \pk_spr_h[20] , \pk_spr_h[13] , \pk_dpr_h[1] , \pk_indx_h[11] , 
        \LDCHK/n3256 , \LBUS/*cell*3982/U31/CONTROL1 , \LBUS/ilt[5] , 
        \SAEXE/n417 , \REGF/RI_SPR[23] , \pk_rwrit_h[25] , \BLU/n1535 , 
        \pk_trba_h[30] , \SADR/pgaddwxyz[13] , rmw12, \CONS/n657 , 
        \pk_indx_h[22] , \SADR/lmtaddr[2] , \pk_rread_h[45] , \LBUS/n_2434 , 
        \REGF/RI_SPR[10] , \pk_trba_h[29] , \pk_indw_h[18] , \pk_idcz_h[1] , 
        \ADOSEL/n4143 , \CODEIF/pgctrinc[4] , \ALUIS/n3641 , \pkbludgh[15] , 
        \CODEIF/n4040 , \pgaluinb[18] , \CODEQ/nqueue1[57] , 
        \REGF/RO_LLPSAS[6] , \LBUS/n1463 , \pk_indy_h[7] , \pk_s6ba_h[2] , 
        \REGF/RO_SRDA[27] , \REGF/RO_SRDA[14] , \REGF/RO_PPCN[11] , 
        \REGF/n8235 , \REGF/n8105 , \REGF/n8095 , \pkdptout[1] , 
        \CODEIF/pfctr[7] , \ALUSHT/pkaluout[27] , \pk_s8ba_h[7] , 
        \REGF/RI_EACC[31] , \REGF/RI_EACC[28] , \REGF/n8122 , \poshtfnc[2] , 
        \CODEQ/nqueue2[27] , \pk_sbba_h[13] , \REGF/RI_PCOL[28] , 
        \REGF/RI_PCOL[31] , pk_ciffh, \REGF/n8212 , ph_shelter_h, 
        \ALUSHT/pkaluout[14] , \LBUS/n1444 , \CODEQ/nqueue2[14] , 
        \CODEIF/n3987 , \pk_rwrit_h[35] , \PDOSEL/n151 , \REGF/n8209 , 
        \pk_dpr_h[8] , \pk_rread_h[55] , \pk_trba_h[20] , \pk_pdo_h[16] , 
        \ALUIS/n3741 , \ph_cpudout[14] , \REGF/RI_SPR[19] , 
        \REGF/pk_s4ba_h[18] , po_trsset_h, \pk_pdo_h[25] , \REGF/n8139 , 
        \pk_trba_h[13] , \pk_indx_h[18] , \REG_2/RETCNT[5] , ph_selldh, 
        \ph_cpudout[27] , \SADR/pgaddwx[20] , \SADR/pgaddwx[13] , 
        \SADR/pgaddyz[6] , \pk_saba_h[6] , \pk_sfba_h[17] , \REGF/RI_PCOH[23] , 
        \REGF/RI_SRA12M[4] , \CONS/SACO[2] , \REGF/RO_PCON[8] , \pk_ada_h[10] , 
        \ph_cpudout[5] , \REGF/RO_PSASL[9] , \pk_ada_h[23] , \BLU/n1582 , 
        \REGF/RI_PCOH[10] , \stream1[10] , \ph_segset_h[7] , 
        \REGF/RI_PCOL[21] , \REGF/RI_EACC[5] , \CODEIF/pfctr[18] , \pgld32[0] , 
        \pgld16[6] , ph_locken_h, \SADR/pgaddxyz[14] , 
        \LBUS/*cell*3982/U185/CONTROL1 , pkalucmf, ph_wrdsrch, \pk_indy_h[15] , 
        \pk_s0ba_h[11] , \REGF/RI_EACC[12] , \LDIS/n3164 , \pk_s9ba_h[17] , 
        \REGF/RI_PCOL[12] , \CODEIF/n3887 , \CODEIF/n3917 , 
        \REGF/pk_indw_h[26] , po_shelter_h1, \REGF/RI_EACC[21] , 
        \CODEQ/nqueue2[37] , \REG_2/ph_retcnt_h[7] , \SADR/pgaddwy[19] , 
        \SADR/pgaddwxz[21] , \SADR/pgaddwxz[12] , \pk_indw_h[22] , 
        \REGF/RO_PPCN[18] , \pgaluinb[22] , ph_d53lth, \pk_indw_h[11] , 
        \pk_s3ba_h[7] , \pk_idcz_h[8] , \REGF/n8195 , \phshtd[4] , 
        \pkdptout[8] , \pgaluinb[11] , \CODEQ/nqueue1[47] , \LDIS/n3143 , 
        \LBUS/srdalth , \CODEIF/n3930 , \BLU/n1509 , \REGF/RI_PCOL[9] , 
        \REGF/RI_TBAI[1] , \BLU/n1499 , \REGF/RO_EST1[1] , \pk_s3ba_h[10] , 
        \ph_segset_h[25] , \stream4[18] , \CODEIF/write_prtect336 , 
        \ALUSHT/pkshtout[20] , \CONS/n535 , \pk_rwrit_h[3] , \REGF/RO_EST2[2] , 
        \pk_pcs2_h[3] , \MAIN/n3620 , ociff, \SADR/pgaddxy[14] , 
        \ph_segset_h[16] , \CONS/n605 , \BLU/n1567 , \REGF/RO_SRDA[9] , 
        \stream4[32] , \ALUSHT/pkshtout[13] , \BLU/n1540 , \pk_pcs2_h[11] , 
        \stream2[0] , \CODEIF/n3979 , \LDIS/ldexcl[14] , \CONS/n622 , 
        \PDOSEL/n79 , \SADR/operand[0] , \pk_sra1_h[22] , \pk_sra1_h[11] , 
        \SADR/pgaddwy[1] , \SADR/pgaddwz[2] , \REGF/RO_PPCN[5] , 
        \pk_idcz_h[14] , \LBUS/*cell*3982/U200/CONTROL1 , \REGF/n8170 , 
        \LDIS/ldexch[16] , \REGF/RI_SRDA[12] , pgperrh, \REGF/RI_DPR[18] , 
        \SADR/m_fadrl[14] , \pgregadrh[2] , \REGF/RI_SRDA[21] , 
        \LDIS/ldexch[25] , \LBUS/n1397 , \LBUS/n1416 , \pk_s9ba_h[9] , 
        \REGF/n8240 , \CODEIF/n3845 , \stream3[40] , \PDOSEL/n103 , 
        \pk_sra1_h[2] , \pk_sra2_h[3] , \stream3[59] , \ADOSEL/n4136 , 
        \CODEIF/n4035 , \ALUIS/n3708 , \ALUIS/n3698 , \LBUS/n1431 , 
        \pk_indx_h[1] , \pk_s2ba_h[0] , \CODEIF/n3862 , \CONS/n739 , 
        \PDOSEL/n124 , \LDCHK/lpex[2] , \REGF/RI_ACC[4] , \CODEIF/n4012 , 
        \REGF/RO_ERRA[6] , \REGF/RI_ACC[19] , \ADOSEL/n4111 , \REGF/n8157 , 
        \pgmuxout[5] , ph_lberr, \CONS/n599 , \pk_seba_h[16] , 
        \REGF/pk_indz_h[25] , \CODEIF/n3971 , ph_exe_dh, seg_config_wr, 
        \CODEQ/nqueue1[11] , \CODEQ/nqueue1[22] , \BLU/n1548 , \pk_indz_h[21] , 
        \SADR/sadr[12] , \pk_sdba_h[15] , \MAIN/sprw_tap2 , \CODEIF/n3956 , 
        \pk_s4ba_h[6] , \pk_psae_h[3] , \REGF/RO_ACC[2] , \PDOSEL/n180 , 
        \LDIS/ldexcl[8] , \pk_idcx_h[6] , \pk_s01l_h[9] , \pk_s45l_h[12] , 
        \LDIS/n3125 , \stream3[25] , \stream3[16] , \SADR/pgaddyz[17] , 
        \pk_indz_h[12] , \SADR/sadr[21] , \pk_s45l_h[21] , \REGF/pk_scti_h[5] , 
        \CODEQ/nqueue2[52] , \pgbluext[30] , \pgbluext[29] , \REGF/n8063 , 
        \MAIN/n3628 , \SADR/pgaddwxy[2] , \SADR/pgaddwxz[1] , 
        \SADR/pgaddxyz[6] , \SADR/pgovfxy , \pk_adb_h[24] , \pk_s2ba_h[13] , 
        \pk_sabl_h[5] , \pgaluinb[3] , \CONS/n591 , \pk_adb_h[17] , 
        \pgaluina[0] , \LBUS/n1439 , \CONS/n731 , \ALUIS/n3727 , 
        \pk_sfba_h[7] , \REGF/RI_PCOH[9] , \pk_rwrit_h[50] , \pk_stdat[19] , 
        \ADOSEL/n4089 , \SAEXE/trsc2_h , \pk_rread_h[30] , \pk_rread_h[29] , 
        \ADOSEL/n4119 , \CONS/n686 , \CONS/n716 , ph_rgfile_h, \BLU/n1474 , 
        \pk_rwrit_h[49] , \REGF/RO_ERRA[15] , \REGF/RO_ERRA[26] , 
        \pk_pcs1_h[2] , \ALUIS/n3700 , \pk_rwrit_h[63] , \ALUIS/n3690 , 
        \REGF/n8178 , ph_initldh, code_area_h, \pgsadrh[4] , \pk_s8ba_h[14] , 
        \REGF/RI_SRA12M[26] , \LDCHK/n3287 , ph_lbussth, \REGF/RO_PCON[28] , 
        \REGF/n8226 , \pk_idcy_h[9] , \ADOSEL/n4150 , \REGF/RO_ACC[16] , 
        \pk_s1ba_h[12] , \ALUSHT/pkshtout[4] , \REGF/RI_SRA12M[15] , 
        \REGF/n8086 , \REGF/n8116 , \pk_s23l_h[31] , \REGF/RO_ACC[25] , 
        \pk_s23l_h[28] , \CODEIF/pgctrinc[10] , \pgsdprlh[9] , 
        \ALUSHT/pkaluout[1] , \REGF/n8131 , \pk_sra2_h[16] , \pk_s5ba_h[1] , 
        \PDOSEL/n142 , \REGF/pk_idcx_h[30] , \REGF/n8201 , \CODEIF/n3994 , 
        \REGF/pk_idcx_h[29] , \PDOSEL/n94 , \pk_rread_h[6] , \ALUIS/n3749 , 
        \LBUS/n1457 , \SADR/segbase[10] , \REGF/RI_SRDA[6] , \pk_pcs1_h[16] , 
        \pk_idcy_h[13] , \ALUIS/n3675 , \pk_s01l_h[27] , \pk_sabl_h[18] , 
        \CODEIF/pfctr415[8] , \CONS/n663 , \CODEIF/n3938 , \BLU/n1501 , 
        \pk_sefl_h[0] , \BLU/n1491 , \SAEXE/n423 , \pk_idcy_h[20] , 
        \LDCHK/n3262 , \SADR/operand[25] , \pk_trba_h[4] , \SADR/pgaddwz[15] , 
        \pk_s01l_h[14] , \REGF/D2_DTFL , \REGF/pk_exco_h[3] , \pk_stdat[1] , 
        \REGF/pk_idcy_h[24] , \pkbludgh[4] , \CONS/n342 , \CONS/n553 , 
        \MAIN/seq_enable , \LDCHK/n3245 , \SADR/pgaddxz[18] , \pgsadrh[22] , 
        \pgsadrh[11] , \REGF/RO_LPSAS2156[1] , \pk_s89l_h[21] , 
        \pk_s89l_h[12] , \pk_idcw_h[17] , ph_saexe_sth, \pgld32[17] , 
        \CONS/n574 , \stream4[57] , \pgld32[24] , \CONS/n644 , \CODEIF/n3904 , 
        \BLU/n1526 , \SADR/operand[16] , \pk_indz_h[6] , \pk_s5ba_h[8] , 
        \CODEIF/n3894 , ph_iyco_h, \ALUIS/n3649 , \CODEIF/pfctr415[14] , 
        \pk_s45l_h[5] , \SADR/operand[9] , \pk_spr_h[4] , \SADR/pgaddxz[22] , 
        \SADR/pgaddwxz[8] , \pk_s0ba_h[4] , \pk_idcx_h[17] , \CONS/n548 , 
        \pk_scba_h[10] , \pk_s23l_h[21] , \pgsdprlh[0] , \REGF/n8186 , 
        ph_tpralt_h, \ALUSHT/pkaluout[8] , \pk_s23l_h[12] , \CODEIF/n3923 , 
        \LDCHK/n3279 , lo_data_lth, \LDIS/n3150 , \REG_2/ncnt2[2] , 
        \pk_idcy_h[0] , \CONS/n678 , \REG_2/ncnt1[1] , \pgsdprlh[12] , 
        \pk_s5ba_h[16] , \pk_saco_lh[3] , \stream4[47] , \ALUIS/n3752 , 
        ret_cont_h, \CONS/n744 , \PDOSEL/n159 , \SADR/pgaddxz[11] , 
        \pk_stdat[8] , \SADR/pgaddwxy[17] , \pgsadrh[18] , \pk_s89l_h[31] , 
        \pgsdprlh[21] , \REGF/RO_LPSAS2156[8] , \pgregadrh[21] , 
        \pgregadrh[12] , \pk_sbba_h[5] , \pk_s89l_h[28] , \pk_sefl_h[9] , 
        \REGF/pk_idcw_h[30] , \REGF/pk_idcw_h[29] , \SADR/lmtaddr[14] , 
        \pk_s67l_h[2] , \pk_s89l_h[3] , \pk_sabl_h[22] , \pk_adb_h[5] , 
        \CODEIF/write_prtect , \MAIN/d_exec_stage , \pk_sabl_h[11] , 
        ph_trslt_h, \REGF/RI_SPR[7] , \CODEIF/pfctr415[1] , \stream3[4] , 
        \pk_dpr_h[17] , \SADR/pgaddwx[5] , ad_latch, \pk_s1ba_h[3] , 
        \pk_s45l_h[31] , \pk_scdl_h[5] , srctype1, \pgaluina[14] , 
        \CODEQ/nqueue2[42] , \pk_s45l_h[28] , \pk_sefl_h[17] , \REGF/n8163 , 
        \pkdptout[16] , ph_timouth, \pgmuxout[24] , \pk_s6ba_h[17] , 
        \ADOSEL/n4125 , \CODEIF/n4026 , \PDOSEL/n110 , \pk_s01l_h[0] , 
        \pk_sefl_h[24] , \pkdptout[25] , \pgmuxout[17] , \LDIS/ldexcl[1] , 
        \CODEIF/n3856 , \REGF/pk_sdba_h[18] , \pgaluina[27] , \LBUS/n1595 , 
        lbus_locken_h, \LBUS/n1405 , \ADOSEL/n4092 , \ADOSEL/n4102 , 
        \CODEQ/nqueue1[32] , \pk_scdl_h[26] , \pk_scdl_h[15] , \pk_idcw_h[2] , 
        \CODEIF/n4001 , \REGF/RI_DPR[2] , \pgbluext[6] , \CODEIF/n3871 , 
        \CONS/SACO[13] , \PDOSEL/n137 , eaccasel, \LBUS/n1422 , 
        \CODEQ/nqueue1[18] , \REGF/n8144 , \REGF/n8078 , \MAIN/n3633 , 
        \pk_scba_h[2] , \pk_s67l_h[14] , \pk_rread_h[13] , \stream2[15] , 
        \CONS/n526 , ph_dec_ch, \REGF/RO_PCON[21] , \pk_s67l_h[27] , 
        \REGF/RI_PCOH[0] , \pk_rwrit_h[40] , \pk_rwrit_h[59] , 
        \pk_rread_h[39] , \pk_rread_h[20] , \stream2[26] , po_reacl_h, 
        \CONS/n616 , \BLU/n1574 , \REGF/RO_PCON[12] , \pk_spr_h[9] , 
        ph_srcadr1_h, \pk_stdat[10] , \LDIS/n3119 , \CONS/n631 , \BLU/n1553 , 
        \SAEXE/sa_start2 , \SADR/pgaddwyz[2] , \pk_s23l_h[7] , 
        \REGF/RO_EACC[3] , \MAIN/n3614 , \LBUS/n1609 , \pgsadrh[15] , 
        \LDCHK/n3230 , \pgaluina[9] , \pgld32[13] , ret_cont_wr, \CONS/n534 , 
        \pk_sbba_h[8] , \pk_s89l_h[25] , \MAIN/n3621 , \pk_stdat[5] , 
        \pk_idcw_h[20] , \REGF/RO_LPSAS2156[5] , \SADR/pgaddwz[22] , 
        \pgsadrh[26] , \pk_s89l_h[16] , \pkbludgh[0] , \BLU/n1566 , 
        \pk_s01l_h[23] , \pk_idcw_h[13] , \stream4[53] , \pgld32[20] , 
        \CONS/n604 , \CODEIF/n3978 , \BLU/n1541 , \SADR/pgaddwz[11] , 
        \SADR/segbase[14] , \pk_idcy_h[17] , \CONS/n623 , \PDOSEL/n78 , 
        \REGF/RI_SRDA[2] , \pk_pcs1_h[12] , \pk_adb_h[8] , \SAEXE/exec_end2 , 
        \pk_s01l_h[10] , \REGF/pk_idcw_h[24] , n10731, \SADR/operand[4] , 
        \stream3[21] , \stream3[12] , \pk_sra2_h[21] , \pk_sefl_h[4] , 
        \pk_s0ba_h[9] , \pk_s45l_h[8] , \REGF/n8171 , \stream3[9] , 
        \pk_sra2_h[12] , \SADR/pgaddwxy[6] , \pk_s5ba_h[5] , \pk_s8ba_h[10] , 
        \pk_rread_h[2] , \ADOSEL/n4137 , \CODEIF/n4034 , \ALUIS/n3699 , 
        ph_exstga_h, \ALUIS/n3709 , \LBUS/n1396 , \LBUS/n1417 , \REGF/n8241 , 
        \CODEIF/n3844 , \REGF/RO_ACC[12] , \PDOSEL/n102 , \ADOSEL/n4110 , 
        \CODEIF/n4013 , \REGF/RI_SRA12M[22] , \LBUS/n1430 , \CONS/n738 , 
        \PDOSEL/n125 , \CODEIF/n3863 , \ALUSHT/pkaluout[5] , 
        \SADR/pgaddwxz[5] , \REGF/RO_ACC[21] , \CODEIF/pgctrinc[14] , 
        \REGF/n8156 , \pgsadrh[0] , \pk_s1ba_h[16] , \REGF/RI_SRA12M[11] , 
        \ALUSHT/pkshtout[0] , \CONS/n598 , \pk_pcs1_h[6] , \ALUIS/n3740 , 
        \pk_dpr_h[30] , \pk_sfba_h[3] , \pk_rwrit_h[54] , \REGF/RO_ERRA[11] , 
        \pk_rread_h[34] , \REGF/n8208 , \pk_dpr_h[29] , \SADR/pgaddyz[20] , 
        \SADR/pgaddyz[13] , \SADR/pgaddxyz[2] , \pk_s67l_h[19] , pk_mpxdh, 
        ph_ebaccwt_h, \REGF/RO_ERRA[22] , \REGF/n8138 , \stream2[18] , 
        \pk_rwrit_h[67] , \pgaluina[4] , \pk_adb_h[20] , \pgaluinb[7] , 
        \pk_s2ba_h[17] , \pk_sabl_h[1] , \pk_indz_h[16] , \SADR/sadr[25] , 
        \SADR/sadr[16] , \pk_s4ba_h[2] , \pk_s45l_h[16] , \pk_adb_h[13] , 
        \BLU/n1583 , \pk_sefl_h[30] , \pk_sefl_h[29] , \LDIS/n3165 , 
        \pk_psae_h[7] , \pk_idcx_h[2] , \REGF/RO_ACC[6] , \pkdptout[31] , 
        \CODEIF/n3886 , \pkdptout[28] , \CODEIF/n3916 , \pk_sdba_h[11] , 
        \pk_s45l_h[25] , \REGF/pk_scti_h[1] , \pgmuxout[29] , \pgmuxout[30] , 
        \pgaluina[19] , \CODEQ/nqueue2[56] , \pk_scdl_h[8] , \pk_sra1_h[6] , 
        \SADR/pgaddwx[8] , \REGF/n8194 , pgpaendp, \CODEQ/nqueue1[15] , 
        \LDIS/n3142 , \pk_sabl_h[8] , \pk_scdl_h[18] , \CODEIF/n3931 , 
        \pk_stdat[14] , \REGF/RO_EACC[7] , \ALUIS/n3667 , \CODEQ/nqueue1[26] , 
        \BLU/n1498 , \BLU/n1508 , pktblcovfh, \BLU/n1483 , \BLU/n1513 , n10736, 
        \SADR/operand[23] , \SADR/operand[21] , \stream3[31] , \stream3[28] , 
        \stream3[0] , \SADR/pgaddwyz[6] , \pk_s23l_h[3] , \LDCHK/n3270 , 
        \LDIS/n3159 , \SAEXE/rf_srcadr1_h , \CONS/n671 , \SAEXE/n431 , 
        ph_d20lth, \pk_scba_h[6] , \pk_adb_h[30] , \CONS/n350 , \CONS/n541 , 
        \pk_adb_h[29] , ph_bit_h, \REGF/RO_PCON[25] , \pk_dpr_h[13] , 
        \pk_s67l_h[10] , \SAEXE/n416 , \pk_rread_h[17] , \stream2[11] , 
        \MAIN/accovf , \LDCHK/n3257 , \CONS/n566 , \pk_spr_h[0] , 
        \pk_dpr_h[20] , \pk_s67l_h[23] , \REGF/RI_PCOH[4] , \REGF/RO_ERRA[18] , 
        \REGF/RO_PCON[16] , \pk_rwrit_h[44] , \BLU/n1534 , \pk_saco_hh[31] , 
        \pk_saco_hh[28] , \CONS/n656 , \pk_trba_h[9] , \SADR/pgaddwx[1] , 
        \pk_scdl_h[11] , \pk_rread_h[24] , \REGF/pk_indz_h[31] , \stream2[22] , 
        \REGF/pk_indz_h[28] , \LBUS/n1462 , \PDOSEL/n177 , \pk_idcw_h[6] , 
        \REGF/RI_DPR[6] , \REGF/n8234 , \pgbluext[2] , \CONS/SACO[17] , 
        \CODEIF/n4041 , \ADOSEL/n4142 , \CODEQ/nqueue1[36] , 
        \SADR/pgaddwz[18] , \SADR/pgaddwxy[20] , \SADR/m_fadrl[6] , 
        \pk_scdl_h[22] , \REGF/n8094 , \REGF/n8104 , \pk_s1ba_h[7] , ph_iwco_h, 
        \pgmuxout[20] , \pk_s6ba_h[13] , \pk_s01l_h[4] , \pk_scdl_h[1] , 
        \pk_sefl_h[13] , \REGF/n8123 , \UPIF/ready_eoc , \pkdptout[12] , 
        \pgaluina[10] , \CODEQ/nqueue2[46] , \pgaluina[23] , \LBUS/n1445 , 
        \pk_sefl_h[20] , \pkdptout[21] , \REGF/n8213 , \pgmuxout[13] , 
        \CODEIF/n3986 , \LDIS/ldexcl[5] , \PDOSEL/n150 , \pk_s01l_h[19] , 
        \pk_s89l_h[7] , \LBUS/ldoe966 , \pk_adb_h[1] , \CONS/n583 , 
        \pk_sabl_h[26] , \SADR/pgaddxz[15] , \SADR/pgaddwxy[13] , 
        \pgregadrh[16] , \SADR/lmtaddr[10] , \pk_sabl_h[15] , \REGF/RI_SPR[3] , 
        \CODEIF/n3878 , \CODEIF/pfctr415[5] , \CONS/n723 , \ALUIS/n3735 , 
        \pk_sbba_h[1] , \pk_s67l_h[6] , \CODEIF/n4008 , \pgsdprlh[16] , 
        ph_trscdech, \pk_saco_lh[7] , \PDOSEL/n119 , \BLU/n1466 , 
        \stream4[43] , \ALUIS/n3682 , \pgld32[29] , \pgld32[30] , \CONS/n704 , 
        \CONS/n694 , \ALUIS/n3712 , rrmw1, \pk_s5ba_h[12] , 
        \REGF/pk_idcy_h[30] , \LDCHK/n3305 , \pkbludgh[9] , \LDCHK/n3295 , 
        \pgsadrh[9] , \pk_scba_h[14] , \REGF/pk_idcy_h[29] , \LDCHK/n3239 , 
        \pk_s23l_h[25] , \pgsdprlh[4] , \REGF/RO_ACC[28] , 
        \MAIN/*cell*4603/U1/CONTROL1 , \REGF/RI_SRA12M[18] , 
        \REGF/RO_PSTA[19] , \ALUSHT/pkshtout[9] , \REGF/n8056 , 
        \pk_s23l_h[16] , \pk_idcx_h[13] , \LBUS/n1600 , \pk_idcy_h[4] , 
        \CONS/n638 , \pk_idcx_h[20] , \CODEIF/pfctr415[10] , \CODEIF/n3963 , 
        \REGF/pk_idcx_h[24] , \LDIS/n3137 , \SADR/operand[12] , 
        \pk_sra2_h[31] , \pk_s0ba_h[0] , sequencial1, \CODEIF/n3944 , 
        \pk_sra2_h[28] , \REGF/n8071 , \pk_spr_h[2] , \SADR/pgaddwxy[22] , 
        \pk_indz_h[2] , \pk_s45l_h[1] , \MAIN/exe_end , \LDCHK/n3292 , 
        \LDCHK/n3302 , \SADR/pgaddwxy[11] , \pgregadrh[14] , 
        \SADR/lmtaddr[12] , \pk_s67l_h[4] , \pk_s89l_h[5] , \pk_sabl_h[24] , 
        \MAIN/ph_rdwr1selh , \pk_adb_h[3] , \REGF/RI_SRDA[9] , \CODEIF/n4028 , 
        \ALUIS/n3715 , \pk_s01l_h[31] , \pk_s01l_h[28] , \ALUIS/n3685 , 
        \REGF/RI_SPR[1] , \CONS/n693 , \CONS/n703 , \pk_sabl_h[17] , 
        \pk_s5ba_h[10] , \pgsdprlh[14] , \CODEIF/n3858 , \CODEIF/pfctr415[7] , 
        \pk_idcw_h[18] , \pk_saco_lh[5] , \REGF/RO_LLPSAS[10] , 
        \LBUS/temp1[2] , \stream4[58] , \stream4[41] , \ALUIS/n3732 , 
        \LBUS/word32odphase , \CONS/n724 , \PDOSEL/n139 , \SADR/pgaddxz[17] , 
        ph_stdatlth, \pk_sbba_h[3] , \pk_scba_h[16] , \pk_s23l_h[27] , 
        \pgsdprlh[6] , \pk_idcx_h[11] , ltffsel, \pgld32[18] , \CONS/n584 , 
        \CONS/n339 , \CONS/n528 , \REGF/n8076 , \pk_s23l_h[14] , 
        \pk_idcx_h[22] , \CODEIF/n3943 , \pk_idcy_h[6] , \LDIS/n3130 , 
        \CONS/n618 , \REGF/RO_ACC[19] , po_wrdsrc_h, \SADR/operand[10] , 
        \pk_sra2_h[19] , \CODEIF/n3964 , \REGF/pk_idcx_h[26] , \LDIS/n3117 , 
        \pk_rread_h[9] , \stream3[33] , \pk_s45l_h[3] , \CODEIF/pfctr415[12] , 
        \LBUS/n1607 , \stream3[19] , \pk_indz_h[0] , ph_trsc_h, \REGF/n8051 , 
        \pk_dpr_h[22] , \pk_dpr_h[11] , \SADR/pgaddyz[18] , \SADR/pgovfwy , 
        \pk_s0ba_h[2] , \pk_stdat[16] , \pk_adb_h[18] , \CONS/n651 , 
        \BLU/n1533 , \SAEXE/bnolth , \REGF/RO_EACC[5] , \ALUIS/n3647 , 
        \SADR/pgaddwyz[4] , \LDCHK/n3250 , \CONS/n561 , \SADR/pgaddxyz[9] , 
        \pk_s23l_h[1] , \SAEXE/n411 , \REGF/n8188 , \CONS/n546 , 
        \pk_scba_h[4] , \pk_s67l_h[12] , \pk_rread_h[15] , \stream2[13] , 
        \MAIN/dprw_inhibith , \LDCHK/n3277 , \REGF/RO_PCON[27] , 
        \pk_rread_h[26] , \stream2[20] , \UPIF/reg_wr , \CONS/n676 , 
        \BLU/n1514 , \SADR/operand[6] , \stream3[2] , \pk_sfba_h[8] , 
        \pk_rwrit_h[46] , \REGF/RO_PCON[14] , \BLU/n1484 , \pk_s67l_h[21] , 
        \REGF/RI_PCOH[6] , \REGF/pk_s2ba_h[18] , \ALUIS/n3660 , \pk_dpr_h[18] , 
        \SADR/pgaddwx[3] , \SADR/m_fadrl[4] , \pk_scdl_h[13] , \pk_idcw_h[4] , 
        \CODEQ/nqueue1[34] , \REGF/RI_DPR[4] , \REGF/n8214 , cif_cont, 
        \CODEIF/n3981 , \CONS/SACO[15] , \PDOSEL/n157 , ph_rmw2h, \LBUS/n1442 , 
        \PDOSEL/n81 , \MAIN/*cell*4603/U15/CONTROL1 , \pk_scdl_h[20] , 
        \REGF/n8124 , \SADR/pgaddxyz[0] , \pk_s1ba_h[5] , \pk_scdl_h[3] , 
        \pk_sefl_h[11] , \pgaluina[12] , \CODEQ/nqueue2[44] , \REGF/n8093 , 
        \REGF/n8103 , \pkdptout[10] , \pk_s4ba_h[9] , \pk_s6ba_h[11] , 
        saenabl2, \pgmuxout[22] , \pgbluext[26] , \pgmuxout[11] , 
        \ADOSEL/n4145 , \LDIS/ldexcl[7] , \pk_sfba_h[1] , \pk_s01l_h[6] , 
        \pkdptout[23] , \REGF/n8233 , \pk_sefl_h[22] , \REGF/RO_ERRA[13] , 
        \pk_idcx_h[9] , \pk_rread_h[36] , \pgaluina[21] , \REGF/n8228 , 
        \BLU/n1584 , \pk_rwrit_h[56] , \pk_s67l_h[31] , \pk_s67l_h[28] , 
        \pk_pcs1_h[4] , \REGF/RO_ERRA[20] , \pk_rwrit_h[65] , \REGF/n8088 , 
        \REGF/n8118 , \SADR/pgaddyz[22] , \SADR/pgaddyz[11] , po_atchk_h, 
        \pk_s23l_h[8] , \pk_adb_h[22] , \pgaluina[6] , \pgaluinb[5] , 
        \pk_adb_h[11] , \LBUS/n1459 , \SADR/sadr[14] , \pk_s2ba_h[15] , 
        \pk_sabl_h[3] , \ALUIS/n3747 , \pk_s4ba_h[0] , \pk_sdba_h[13] , 
        \pk_s45l_h[14] , \pk_psae_h[5] , \pk_idcx_h[0] , \REGF/RO_ACC[4] , 
        \pgmuxout[18] , \CODEIF/n3936 , \pgaluina[28] , \pgaluina[31] , 
        \LDIS/n3145 , ph_ldaoutenh1, \pk_sra1_h[4] , \pk_indz_h[14] , 
        \pk_s45l_h[27] , \pk_sefl_h[18] , \SADR/sadr[27] , \REGF/pk_scti_h[3] , 
        \CODEQ/nqueue2[54] , \REGF/n8193 , \pkdptout[19] , \pk_scdl_h[30] , 
        \pk_scdl_h[29] , \CODEQ/nqueue1[17] , \REGF/RO_TRCO[26] , 
        \pgbluext[9] , \CODEIF/n3911 , ph_exe_bh, \CODEQ/nqueue1[24] , 
        \BLU/n1528 , \CODEIF/n3881 , \LDIS/n3162 , \SADR/pgaddwz[20] , 
        \SADR/pgaddwxy[18] , \pgsadrh[24] , \pgsadrh[17] , \pk_s89l_h[27] , 
        \pk_stdat[7] , \pk_idcw_h[22] , \pkbludgh[2] , \REGF/RO_LPSAS2156[7] , 
        \pk_idcw_h[11] , \pgld32[11] , \stream4[51] , \stream4[48] , 
        \pgld32[22] , \CONS/n624 , \SADR/segbase[16] , \pk_s89l_h[14] , 
        \BLU/n1546 , \REGF/RI_SRDA[0] , \MAIN/ADROVH , \pk_pcs1_h[10] , 
        \UPIF/tr_count_lt , \pk_idcy_h[15] , \CODEIF/n3958 , \CONS/n603 , 
        \pk_s01l_h[21] , \REGF/RI_SPR[8] , \pk_sefl_h[6] , \BLU/n1561 , 
        \SADR/operand[27] , \SADR/operand[19] , \SADR/pgaddwz[13] , 
        \pk_s01l_h[12] , \REGF/pk_idcw_h[26] , up_data_lth, ph_dregsl_h, 
        \MAIN/c_exec_stage , \MAIN/n3626 , \CONS/n533 , \stream3[23] , 
        \stream3[10] , \pk_indz_h[9] , \REGF/n8151 , \pk_sra2_h[23] , 
        \pk_sra2_h[10] , \pk_s5ba_h[7] , \CODEIF/n3864 , \PDOSEL/n122 , 
        \MAIN/excep_valid , \LBUS/n1437 , \pk_rread_h[0] , \CODEIF/n4014 , 
        \ADOSEL/n4087 , \ALUIS/n3729 , \ADOSEL/n4117 , \stream3[6] , 
        \pk_dpr_h[15] , \pk_sra1_h[9] , \SADR/pgaddwxy[4] , \SADR/pgaddwxz[7] , 
        \pgsadrh[2] , \pk_s8ba_h[12] , \REGF/RI_SRA12M[20] , 
        \REGF/RO_PSTA[21] , \CODEIF/n3843 , \PDOSEL/n105 , \LBUS/n1410 , 
        \LBUS/n1391 , \CONS/n688 , \CONS/n718 , \ADOSEL/n4130 , 
        \REGF/RO_ACC[10] , \ph_pdis_h[10] , \CODEIF/n4033 , phadrinch, 
        \pk_s1ba_h[14] , \pk_idcx_h[18] , \ALUSHT/pkshtout[2] , 
        \REGF/RI_SRA12M[13] , \REGF/n8176 , \REGF/RO_ACC[23] , 
        \CODEIF/pgctrinc[16] , \pk_indz_h[19] , \pk_s1ba_h[1] , \LDCHK/n3289 , 
        \ALUSHT/pkaluout[7] , \pk_sefl_h[15] , \REGF/n8143 , \pgmuxout[26] , 
        \pkdptout[14] , \SADR/sadr[19] , \pk_s01l_h[2] , \pk_scdl_h[7] , 
        \pgaluina[16] , \CODEQ/nqueue2[40] , \CODEQ/nqueue2[59] , 
        \pk_sefl_h[26] , \pgaluina[25] , \CMPX/n1048 , \LBUS/n1425 , 
        \pk_s45l_h[19] , \pkdptout[27] , \pk_s6ba_h[15] , \CODEIF/n3876 , 
        \REGF/RO_ACC[9] , \pgmuxout[15] , \PDOSEL/n130 , \LDIS/ldexcl[3] , 
        \ADOSEL/n4095 , \ADOSEL/n4105 , \CODEIF/n4006 , \SADR/pgaddwx[7] , 
        \pk_scdl_h[17] , \LBUS/n1402 , \LBUS/n1592 , \PDOSEL/n117 , 
        \BLU/n1468 , \pk_idcw_h[0] , pk_sign_h, \pgbluext[4] , \CONS/SACO[11] , 
        \REGF/RI_DPR[0] , \CODEIF/n3851 , \ADOSEL/n4122 , \CODEIF/n4021 , 
        \CODEQ/nqueue1[29] , \CODEQ/nqueue1[30] , \pk_scba_h[0] , 
        \pk_scdl_h[24] , \REGF/n8164 , \REGF/RO_PCON[23] , \pk_s67l_h[16] , 
        ph_schvx_h, \LDCHK/n3237 , ph_dec_ah, \UPIF/n1046 , \pk_rread_h[11] , 
        step3_cf, \pk_rwrit_h[68] , \REGF/n8058 , \MAIN/n3613 , 
        \SADR/pgaddwyz[0] , \pk_s67l_h[25] , \pk_pcs1_h[9] , \REGF/RI_PCOH[2] , 
        \pk_rwrit_h[42] , \REGF/RO_PCON[10] , \BLU/n1554 , \pk_stdat[12] , 
        \pk_rread_h[22] , \MAIN/dec_end , \CONS/n636 , \REGF/RO_EACC[1] , 
        \LDIS/n3139 , \BLU/n1573 , \CONS/n611 , \pk_s23l_h[5] , 
        \CODEIF/pfctr415[16] , \pgaluinb[8] , \MAIN/n3634 , \CONS/n521 , 
        \ALUIS/n3669 , \LDIS/n3157 , \CODEIF/n3924 , \SADR/operand[14] , 
        \pk_indz_h[4] , \pk_s0ba_h[6] , po_mode01_h, \REGF/n8181 , 
        \SAEXE/*cell*3651/U11/CONTROL1 , \pk_spr_h[6] , \SADR/pgaddxz[20] , 
        \SADR/pgaddwxy[9] , \pk_scba_h[12] , \pk_s45l_h[7] , \pk_saseo_h[1] , 
        \LDCHK/n3259 , \SAEXE/n418 , \pk_s23l_h[23] , \pk_s23l_h[10] , 
        \pgsdprlh[2] , \pk_idcx_h[15] , \CONS/n568 , \pk_s89l_h[19] , 
        \pk_idcy_h[2] , \CONS/n658 , \REG_2/ncnt2[0] , \CODEIF/n3893 , 
        \CODEIF/n3903 , \PDOSEL/n179 , \pk_saco_lh[1] , \REGF/RO_LLPSAS[14] , 
        \stream4[45] , \REG_2/n435 , \SADR/pgaddxz[13] , \pk_sbba_h[7] , 
        \pgsdprlh[10] , \pgsdprlh[23] , \pk_s5ba_h[14] , \pgregadrh[10] , 
        \pk_s89l_h[1] , \pk_sabl_h[20] , \pk_adb_h[7] , ph_d76lth, 
        \RSTGN/CRST_2H , \stream3[27] , \stream3[14] , \SADR/pgaddwxy[15] , 
        \pgregadrh[23] , wacc, \CODEIF/pfctr415[3] , \CODEIF/n3988 , 
        \SADR/pgaddwxy[0] , \pk_s8ba_h[16] , \pk_s23l_h[19] , \pk_s67l_h[0] , 
        \pk_sabl_h[13] , \REGF/RI_SPR[5] , \CONS/n743 , \pk_idcy_h[18] , 
        \LDCHK/pchkenh , \REGF/RO_ACC[14] , ph_adrwtenh, \LBUS/n1450 , 
        \REGF/RI_SRA12M[24] , \PDOSEL/n145 , \REGF/n8206 , \CODEIF/n3993 , 
        \pgfdout[0] , \ALUSHT/pkaluout[3] , \SADR/pgaddwxz[3] , 
        \REGF/RI_SRA12M[17] , \REGF/RO_ACC[27] , \CODEIF/pgctrinc[12] , 
        \REGF/RO_PSTA[16] , \pgsadrh[6] , \pk_s1ba_h[10] , \REGF/n8136 , 
        \ALUSHT/pkshtout[6] , \REGF/n8081 , \REGF/n8111 , \pk_sra2_h[14] , 
        \SADR/pgaddwz[17] , \SADR/segbase[12] , \pk_s5ba_h[3] , 
        \pk_s01l_h[25] , \pk_rread_h[4] , \ADOSEL/n4157 , \REGF/n8221 , 
        pkaluovf, \PDOSEL/n162 , \BLU/n1521 , \CODEIF/n3888 , \CODEIF/n3918 , 
        \CONS/n643 , \pk_s67l_h[9] , \pk_pcs1_h[14] , \pk_idcy_h[11] , 
        \ALUIS/n3655 , \pk_s89l_h[8] , \REGF/RI_SRDA[4] , \CONS/n573 , 
        \pgregadrh[19] , \pk_s01l_h[16] , \pk_sabl_h[29] , \REGF/pk_exco_h[1] , 
        \pk_sabl_h[30] , \ALUSHT/slaovf , pk_pcon31_h, \SADR/operand[2] , 
        \pk_sra1_h[0] , \pk_trba_h[6] , \pgsadrh[13] , \pk_s89l_h[23] , 
        \pk_sefl_h[2] , \pk_idcy_h[22] , \pgld32[15] , \LDCHK/n3242 , 
        \CONS/n554 , \CONS/n345 , \pgsadrh[20] , \pk_stdat[3] , 
        \REGF/pk_idcy_h[26] , \REGF/RO_LPSAS2156[3] , \pkbludgh[6] , 
        \LDCHK/n3265 , \pk_saco_lh[8] , cnt_write_h, \SAEXE/n424 , \BLU/n1496 , 
        \BLU/n1506 , \SADR/m_fadrl[9] , \pk_s89l_h[10] , \pgsdprlh[19] , 
        \stream4[55] , rmw21, \pgld32[26] , \CONS/n664 , \ALUIS/n3672 , 
        \pk_idcw_h[15] , \REGF/n8064 , \LBUS/n1632 , \LDIS/n3122 , 
        \CODEQ/nqueue1[13] , \pk_indz_h[23] , \pk_idcw_h[9] , 
        \REGF/pk_indz_h[27] , \REGF/pk_s6ba_h[18] , \CODEIF/n3951 , 
        \CONS/SACO[18] , \REGF/RI_DPR[9] , ph_wdstenh, \BLU/n1568 , 
        \CODEQ/nqueue1[39] , \CODEQ/nqueue1[20] , srcbsel, \pk_indz_h[10] , 
        \SADR/sadr[23] , \SADR/sadr[10] , \pk_s45l_h[10] , \pk_psae_h[1] , 
        \pk_idcx_h[4] , \PDOSEL/n76 , \REGF/RO_ACC[0] , \pk_s4ba_h[4] , 
        \CODEIF/n3976 , \pk_sdba_h[17] , \ALUSHT/n3112 , \pk_s1ba_h[8] , 
        \REGF/pk_scti_h[7] , \CODEQ/nqueue2[50] , \CODEQ/nqueue2[49] , 
        \pk_s45l_h[23] , \MAIN/*cell*4603/U7/CONTROL1 , \SADR/pgaddyz[15] , 
        \SADR/pgaddwyz[9] , \LDCHK/n3280 , \LDCHK/n3310 , \pk_adb_h[26] , 
        \pgaluina[2] , \pgaluinb[1] , \SAEXE/adovflth2 , \SADR/pgaddxyz[4] , 
        \pk_s2ba_h[11] , \REGF/RO_EACC[8] , \ADOSEL/n4139 , \ALUIS/n3697 , 
        \ALUIS/n3707 , \pk_scba_h[9] , \pk_sfba_h[5] , \pk_sabl_h[7] , accasel, 
        \pk_pcs1_h[0] , \pk_adb_h[15] , \LBUS/n1419 , \LBUS/n1398 , 
        \BLU/n1473 , \CONS/n711 , \CONS/n681 , \ALUIS/n3720 , 
        \REGF/RO_PCON[19] , \pk_rwrit_h[52] , \REGF/RO_ERRA[17] , 
        \pk_rread_h[32] , ph_sprsel2_h, \UPIF/write_by_h , \CONS/n736 , 
        \CONS/n596 , \REGF/RO_ERRA[24] , \pk_rread_h[18] , \pk_rwrit_h[61] , 
        \REGF/n8158 , \MCD/insdec_1/n4197 , \MCD/insdec_1/n4169 , 
        \MCD/insdec_1/n4185 , \MCD/insdec_1/n4160 , \MCD/insdec_1/n4277 , 
        \MCD/insdec_1/n4250 , \MCD/insdec_1/n4202 , \MCD/insdec_1/n4219 , 
        \MCD/insdec_1/n4225 , \MCD/insdec_1/n4259 , \MCD/insdec_1/n4237 , 
        \MCD/insdec_1/n4210 , \MCD/insdec_1/n4280 , \MCD/insdec_1/n4172 , 
        \MCD/insdec_1/n4265 , \MCD/insdec_1/n4245 , \MCD/insdec_1/n4242 , 
        \MCD/insdec_1/n4175 , \MCD/insdec_1/n4262 , \MCD/insdec_1/n4190 , 
        \MCD/insdec_1/n4217 , \MCD/insdec_1/n4230 , \MCD/insdec_1/n4279 , 
        \MCD/insdec_1/n4196 , \MCD/insdec_1/n4167 , \MCD/insdec_1/n4182 , 
        \MCD/insdec_1/n4199 , \MCD/insdec_1/n4205 , \MCD/insdec_1/n4222 , 
        \MCD/insdec_1/n4239 , \MCD/insdec_1/n4257 , \MCD/insdec_1/n4161 , 
        \MCD/insdec_1/n4184 , \MCD/insdec_1/n4223 , \MCD/insdec_1/n4191 , 
        \MCD/insdec_1/ciff , \MCD/insdec_1/n4270 , \MCD/insdec_1/n4278 , 
        \MCD/insdec_1/n4216 , \MCD/insdec_1/n4231 , \MCD/insdec_1/n4166 , 
        \MCD/insdec_1/n4174 , \MCD/insdec_1/n4244 , \MCD/insdec_1/n4256 , 
        \MCD/insdec_1/n4263 , \MCD/insdec_1/n4183 , \MCD/insdec_1/n4271 , 
        \MCD/insdec_1/n4238 , \MCD/insdec_1/n4198 , \MCD/insdec_1/n4204 , 
        \MCD/insdec_1/n4203 , \MCD/insdec_1/n4224 , \MCD/insdec_1/n4218 , 
        \MCD/insdec_1/n4276 , \MCD/insdec_1/n4251 , \MCD/insdec_1/n4173 , 
        \MCD/insdec_1/n4264 , \MCD/insdec_1/n4243 , \MCD/insdec_1/n4195 , 
        \MCD/insdec_1/n4171 , \MCD/insdec_1/n4168 , \MCD/insdec_1/bacc , 
        \MCD/insdec_1/n4281 , \MCD/insdec_1/n4211 , \MCD/insdec_1/n4236 , 
        \MCD/insdec_1/n4258 , \MCD/insdec_1/n4213 , \MCD/insdec_1/n4163 , 
        \MCD/insdec_1/n4186 , \MCD/insdec_1/n4253 , \MCD/insdec_1/n4274 , 
        \MCD/insdec_1/n4178 , \MCD/insdec_1/n4201 , \MCD/insdec_1/n4226 , 
        \MCD/insdec_1/n4248 , \MCD/insdec_1/n4234 , \MCD/insdec_1/n4194 , 
        \MCD/insdec_1/n4208 , \MCD/insdec_1/n4241 , \MCD/insdec_1/n4158 , 
        \MCD/insdec_1/n4176 , \MCD/insdec_1/n4266 , \MCD/insdec_1/n4246 , 
        \MCD/insdec_1/n4261 , \MCD/insdec_1/n4188 , \MCD/insdec_1/n4193 , 
        \MCD/insdec_1/n4214 , \MCD/insdec_1/n4228 , \MCD/insdec_1/n4233 , 
        \MCD/insdec_1/n4268 , \MCD/insdec_1/n4181 , \MCD/insdec_1/n4206 , 
        \MCD/insdec_1/n4221 , \MCD/insdec_1/n4164 , \MCD/insdec_1/n4254 , 
        \MCD/insdec_1/n4273 , \MCD/insdec_1/n4189 , \MCD/insdec_1/n4215 , 
        \MCD/insdec_1/n4232 , \MCD/insdec_1/n4165 , \MCD/insdec_1/n4177 , 
        \MCD/insdec_1/n4192 , \MCD/insdec_1/n4229 , \MCD/insdec_1/n4247 , 
        \MCD/insdec_1/n4260 , \MCD/insdec_1/n4255 , \MCD/insdec_1/n4272 , 
        \MCD/insdec_1/n4159 , \MCD/insdec_1/n4180 , \MCD/insdec_1/n4207 , 
        \MCD/insdec_1/n4220 , \MCD/insdec_1/n4269 , \MCD/insdec_1/n4179 , 
        \MCD/insdec_1/n4249 , \MCD/insdec_1/n4200 , \MCD/insdec_1/n4227 , 
        \MCD/insdec_1/n4162 , \MCD/insdec_1/n4187 , \MCD/insdec_1/n4170 , 
        \MCD/insdec_1/n4252 , \MCD/insdec_1/n4275 , \MCD/insdec_1/n4240 , 
        \MCD/insdec_1/n4267 , \MCD/insdec_1/n4282 , \MCD/insdec_1/n4209 , 
        \MCD/insdec_1/n4212 , \MCD/insdec_1/n4235 , \MAIN/MCD/nst[0] , 
        \MAIN/MCD/n3368 , \MAIN/MCD/n3373 , \MAIN/MCD/dst[0] , 
        \MAIN/MCD/n3396 , \MAIN/MCD/n3384 , \MAIN/MCD/n3367 , 
        \MAIN/MCD/dst[2] , \MAIN/MCD/n3383 , \MAIN/MCD/n3391 , 
        \MAIN/MCD/n3398 , \MAIN/MCD/n3374 , \MAIN/MCD/n3382 , \MAIN/MCD/n3369 , 
        \MAIN/MCD/n3375 , \MAIN/MCD/n3390 , \MAIN/MCD/nst[1] , 
        \MAIN/MCD/n3372 , \MAIN/MCD/n3397 , \MAIN/MCD/n3370 , \MAIN/MCD/n3385 , 
        \MAIN/MCD/dst[1] , \MAIN/MCD/nst[2] , \MAIN/MCD/n3379 , 
        \MAIN/MCD/n3395 , \MAIN/MCD/n3380 , \MAIN/MCD/n3387 , \MAIN/MCD/n3389 , 
        \MAIN/MCD/n3371 , \MAIN/MCD/n3376 , \MAIN/MCD/n3377 , \MAIN/MCD/n3392 , 
        \MAIN/MCD/n3381 , \MAIN/MCD/n3388 , \MAIN/MCD/n3393 , \MAIN/MCD/n3394 , 
        \MAIN/MCD/stage_a154 , \MAIN/MCD/n3386 , \MAIN/MCD/n3378 , 
        \REGF/pbmemcnt1/n6441 , \REGF/pbmemcnt1/upcnt_data283[6] , 
        \REGF/pbmemcnt1/down_data274[2] , \REGF/pbmemcnt1/down_data[5] , 
        \REGF/pbmemcnt1/upcnt_data283[2] , \REGF/pbmemcnt1/time_delay400 , 
        \REGF/pbmemcnt1/n6445 , \REGF/pbmemcnt1/n6495 , 
        \REGF/pbmemcnt1/upcnt_data[3] , \REGF/pbmemcnt1/down_data274[6] , 
        \REGF/pbmemcnt1/down_data[1] , \REGF/pbmemcnt1/upcnt_data[7] , 
        \REGF/pbmemcnt1/upcnt_data283[0] , \REGF/pbmemcnt1/upcnt_data[5] , 
        \REGF/pbmemcnt1/upcnt_data392[11] , \REGF/pbmemcnt1/n6442 , 
        \REGF/pbmemcnt1/down_data274[4] , \REGF/pbmemcnt1/upcnt_data283[9] , 
        \REGF/pbmemcnt1/down_data[3] , \REGF/pbmemcnt1/n401 , 
        \REGF/pbmemcnt1/upcnt_data[1] , \REGF/pbmemcnt1/n6443 , 
        \REGF/pbmemcnt1/upcnt_data283[10] , \REGF/pbmemcnt1/upcnt_data283[4] , 
        \REGF/pbmemcnt1/n6450 , \REGF/pbmemcnt1/down_data[7] , 
        \REGF/pbmemcnt1/upcnt_data392[5] , \REGF/pbmemcnt1/down_data274[0] , 
        \REGF/pbmemcnt1/upcnt_data[8] , \REGF/pbmemcnt1/down_data404[3] , 
        \REGF/pbmemcnt1/upcnt_data392[8] , \REGF/pbmemcnt1/upcnt_data392[1] , 
        \REGF/pbmemcnt1/n6451 , \REGF/pbmemcnt1/upcnt_data[11] , 
        \REGF/pbmemcnt1/down_data404[7] , \REGF/pbmemcnt1/end_flag , 
        \REGF/pbmemcnt1/down_data404[5] , \REGF/pbmemcnt1/n6494 , 
        \REGF/pbmemcnt1/upcnt_data392[3] , \REGF/pbmemcnt1/upcnt_data392[7] , 
        \REGF/pbmemcnt1/down_data404[1] , \REGF/pbmemcnt1/n6444 , 
        \REGF/pbmemcnt1/n393[0] , \REGF/pbmemcnt1/upcnt_data392[6] , 
        \REGF/pbmemcnt1/down_data404[0] , \REGF/pbmemcnt1/down_data404[4] , 
        \REGF/pbmemcnt1/upcnt_data392[2] , \REGF/pbmemcnt1/n6446 , 
        \REGF/pbmemcnt1/upcnt_data392[0] , \REGF/pbmemcnt1/upcnt_data[10] , 
        \REGF/pbmemcnt1/n6447 , \REGF/pbmemcnt1/down_data404[6] , 
        \REGF/pbmemcnt1/upcnt_data392[9] , \REGF/pbmemcnt1/upcnt_data392[4] , 
        \REGF/pbmemcnt1/n6453 , \REGF/pbmemcnt1/upcnt_data283[11] , 
        \REGF/pbmemcnt1/upcnt_data392[10] , \REGF/pbmemcnt1/n6448 , 
        \REGF/pbmemcnt1/down_data404[2] , \REGF/pbmemcnt1/upcnt_data283[5] , 
        \REGF/pbmemcnt1/upcnt_data[0] , \REGF/pbmemcnt1/down_data[6] , 
        \REGF/pbmemcnt1/upcnt_data283[8] , \REGF/pbmemcnt1/upcnt_data283[1] , 
        \REGF/pbmemcnt1/upcnt_data[9] , \REGF/pbmemcnt1/down_data274[1] , 
        \REGF/pbmemcnt1/upcnt_data[4] , \REGF/pbmemcnt1/n6449 , 
        \REGF/pbmemcnt1/n6452 , \REGF/pbmemcnt1/down_data274[5] , 
        \REGF/pbmemcnt1/down_data[2] , \REGF/pbmemcnt1/upcnt_data283[7] , 
        \REGF/pbmemcnt1/upcnt_data283[3] , \REGF/pbmemcnt1/n405[0] , 
        \REGF/pbmemcnt1/upcnt_data[6] , \REGF/pbmemcnt1/down_data274[7] , 
        \REGF/pbmemcnt1/down_data[0] , \REGF/pbmemcnt1/down_data274[3] , 
        \REGF/pbmemcnt1/down_data[4] , \REGF/pbmemcnt1/upcnt_data[2] , 
        \SAEXE/SRCWT/nwst[1] , \SAEXE/SRCWT/ewst[0] , \SAEXE/SRCWT/n85 , 
        \SAEXE/SRCWT/nwst[0] , \MCD/adsel_1/n4292 , \MCD/adsel_1/n4302 , 
        \MCD/adsel_1/n4325 , \MCD/adsel_1/n4289 , \MCD/adsel_1/n4319 , 
        \MCD/adsel_1/n4310 , \MCD/adsel_1/n4350 , \MCD/adsel_1/n4342 , 
        \MCD/adsel_1/n4365 , \MCD/adsel_1/n4337 , \MCD/adsel_1/n4359 , 
        \MCD/adsel_1/n4283 , \MCD/adsel_1/n4287 , \MCD/adsel_1/n4317 , 
        \MCD/adsel_1/n4330 , \MCD/adsel_1/n4286 , \MCD/adsel_1/n4295 , 
        \MCD/adsel_1/n4345 , \MCD/adsel_1/n4362 , \MCD/adsel_1/n4357 , 
        \MCD/adsel_1/n4339 , \MCD/adsel_1/n4305 , \MCD/adsel_1/n4322 , 
        \MCD/adsel_1/n4363 , \MCD/adsel_1/ciff , \MCD/adsel_1/n4344 , 
        \MCD/adsel_1/n4288 , \MCD/adsel_1/n4294 , \MCD/adsel_1/n4304 , 
        \MCD/adsel_1/n4316 , \MCD/adsel_1/n4331 , \MCD/adsel_1/n4323 , 
        \MCD/adsel_1/n4338 , \MCD/adsel_1/n4351 , \MCD/adsel_1/n4356 , 
        \MCD/adsel_1/n4291 , \MCD/adsel_1/n4293 , \MCD/adsel_1/n4318 , 
        \MCD/adsel_1/n4324 , \MCD/adsel_1/n4303 , \MCD/adsel_1/n4311 , 
        \MCD/adsel_1/n4336 , \MCD/adsel_1/n4358 , \MCD/adsel_1/bacc , 
        \MCD/adsel_1/n4343 , \MCD/adsel_1/n4348 , \MCD/adsel_1/n4364 , 
        \MCD/adsel_1/n4301 , \MCD/adsel_1/n4326 , \MCD/adsel_1/n4353 , 
        \MCD/adsel_1/n4366 , \MCD/adsel_1/n4341 , \MCD/adsel_1/n4298 , 
        \MCD/adsel_1/n4308 , \MCD/adsel_1/n4313 , \MCD/adsel_1/n4334 , 
        \MCD/adsel_1/n4284 , \MCD/adsel_1/n4333 , \MCD/adsel_1/n4285 , 
        \MCD/adsel_1/n4296 , \MCD/adsel_1/n4314 , \MCD/adsel_1/n4328 , 
        \MCD/adsel_1/n4346 , \MCD/adsel_1/n4354 , \MCD/adsel_1/n4361 , 
        \MCD/adsel_1/n4306 , \MCD/adsel_1/n4321 , \MCD/adsel_1/n4347 , 
        \MCD/adsel_1/n4360 , \MCD/adsel_1/n4315 , \MCD/adsel_1/n4329 , 
        \MCD/adsel_1/n4332 , \MCD/adsel_1/n4297 , \MCD/adsel_1/n4320 , 
        \MCD/adsel_1/n4307 , \MCD/adsel_1/n4355 , \MCD/adsel_1/n4352 , 
        \MCD/adsel_1/n4290 , \MCD/adsel_1/n4300 , \MCD/adsel_1/n4299 , 
        \MCD/adsel_1/n4312 , \MCD/adsel_1/n4327 , \MCD/adsel_1/n4349 , 
        \MCD/adsel_1/n4335 , \MCD/adsel_1/n4309 , \MCD/adsel_1/n4340 , 
        \LBUS/phsdlt_1/nrt[2] , \LBUS/phsdlt_1/n1012 , \LBUS/phsdlt_1/n1015 , 
        \LBUS/phsdlt_1/n1013 , \LBUS/phsdlt_1/nrt[0] , \LBUS/phsdlt_1/n1014 , 
        \LBUS/phsdlt_1/nrt[1] , \CONS/phsegsel_1/n328 , \CONS/phsegsel_1/n330 , 
        \CONS/phsegsel_1/n336 , \CONS/phsegsel_1/n337 , \CONS/phsegsel_1/n331 , 
        \CONS/phsegsel_1/n333 , \CONS/phsegsel_1/n329 , \CONS/phsegsel_1/n334 , 
        \CONS/phsegsel_1/n335 , \CONS/phsegsel_1/n332 , 
        \REG_2/SATIME/count97[20] , \REG_2/SATIME/count97[16] , 
        \REG_2/SATIME/count[2] , \REG_2/SATIME/count[17] , \REG_2/SATIME/n245 , 
        \REG_2/SATIME/n262 , \REG_2/SATIME/count97[12] , \REG_2/SATIME/n230 , 
        \REG_2/SATIME/count[6] , \REG_2/SATIME/count[20] , 
        \REG_2/SATIME/count[13] , \REG_2/SATIME/n257 , \REG_2/SATIME/n270 , 
        \REG_2/SATIME/n239 , \REG_2/SATIME/count97[19] , 
        \REG_2/SATIME/count[18] , \REG_2/SATIME/n250 , \REG_2/SATIME/n277 , 
        \REG_2/SATIME/dda0 , \REG_2/SATIME/count97[10] , 
        \REG_2/SATIME/count[11] , \REG_2/SATIME/count[4] , \REG_2/SATIME/n237 , 
        \REG_2/SATIME/n259 , \REG_2/SATIME/count[9] , 
        \REG_2/SATIME/count97[14] , \REG_2/SATIME/n242 , 
        \REG_2/SATIME/count[15] , \REG_2/SATIME/count[0] , \REG_2/SATIME/n265 , 
        \REG_2/SATIME/n227 , \REG_2/SATIME/count145[20] , 
        \REG_2/SATIME/count145[18] , \REG_2/SATIME/count145[15] , 
        \REG_2/SATIME/count97[7] , \REG_2/SATIME/count145[0] , 
        \REG_2/SATIME/n251 , \REG_2/SATIME/n276 , \REG_2/SATIME/count145[9] , 
        \REG_2/SATIME/dda1 , \REG_2/SATIME/count145[13] , 
        \REG_2/SATIME/count145[11] , \REG_2/SATIME/count145[4] , 
        \REG_2/SATIME/count97[3] , \REG_2/SATIME/n243 , \REG_2/SATIME/n264 , 
        \REG_2/SATIME/n258 , \REG_2/SATIME/count97[8] , \REG_2/SATIME/n236 , 
        \REG_2/SATIME/n228 , \REG_2/SATIME/count145[17] , 
        \REG_2/SATIME/count145[6] , \REG_2/SATIME/n231 , 
        \REG_2/SATIME/count97[1] , \REG_2/SATIME/n244 , \REG_2/SATIME/n263 , 
        \REG_2/SATIME/n238 , \REG_2/SATIME/n256 , \REG_2/SATIME/n271 , 
        \REG_2/SATIME/count97[5] , \REG_2/SATIME/count145[2] , 
        \REG_2/SATIME/count145[19] , \REG_2/SATIME/count145[16] , 
        \REG_2/SATIME/ph_timouth117 , \REG_2/SATIME/n261 , \REG_2/SATIME/n246 , 
        \REG_2/SATIME/count145[12] , \REG_2/SATIME/count97[4] , 
        \REG_2/SATIME/count145[3] , \REG_2/SATIME/n233 , 
        \REG_2/SATIME/count97[9] , \REG_2/SATIME/count145[7] , 
        \REG_2/SATIME/n268 , \REG_2/SATIME/count97[2] , 
        \REG_2/SATIME/count97[0] , \REG_2/SATIME/n254 , \REG_2/SATIME/n273 , 
        \REG_2/SATIME/count145[14] , \REG_2/SATIME/count145[10] , 
        \REG_2/SATIME/count145[5] , \REG_2/SATIME/n248 , \REG_2/SATIME/n253 , 
        \REG_2/SATIME/n274 , \REG_2/SATIME/count97[6] , 
        \REG_2/SATIME/count145[1] , \REG_2/SATIME/n234 , \REG_2/SATIME/n241 , 
        \REG_2/SATIME/n266 , \REG_2/SATIME/count145[8] , \REG_2/SATIME/n249 , 
        \REG_2/SATIME/count[8] , \REG_2/SATIME/count97[15] , 
        \REG_2/SATIME/count[1] , \REG_2/SATIME/count[14] , \REG_2/SATIME/dda2 , 
        \REG_2/SATIME/n252 , \REG_2/SATIME/n275 , \REG_2/SATIME/count97[18] , 
        \REG_2/SATIME/count[19] , \REG_2/SATIME/n240 , \REG_2/SATIME/n267 , 
        \REG_2/SATIME/count97[11] , \REG_2/SATIME/n235 , \REG_2/SATIME/n232 , 
        \REG_2/SATIME/count[5] , \REG_2/SATIME/count[10] , 
        \REG_2/SATIME/count97[13] , \REG_2/SATIME/count[7] , 
        \REG_2/SATIME/count[12] , \REG_2/SATIME/n247 , \REG_2/SATIME/n260 , 
        \REG_2/SATIME/n229 , \REG_2/SATIME/count97[17] , 
        \REG_2/SATIME/count[3] , \REG_2/SATIME/count[16] , \REG_2/SATIME/n255 , 
        \REG_2/SATIME/n272 , \REG_2/SATIME/n269 , \SAEXE/RFIO/cnt4out[3] , 
        \SAEXE/RFIO/cnt4out[2] , \SAEXE/RFIO/cnt4out[0] , \SAEXE/RFIO/reloadh , 
        \SAEXE/RFIO/nfst[2] , \SAEXE/RFIO/phadrovfh , \SAEXE/RFIO/n379 , 
        \SAEXE/RFIO/n362 , \SAEXE/RFIO/n387 , \SAEXE/RFIO/n406 , 
        \SAEXE/RFIO/n395 , \SAEXE/RFIO/n357 , \SAEXE/RFIO/n370 , 
        \SAEXE/RFIO/n389 , \SAEXE/RFIO/*cell*3735/U62/CONTROL2 , 
        \SAEXE/RFIO/n408 , \SAEXE/RFIO/n377 , \SAEXE/RFIO/n392 , 
        \SAEXE/RFIO/cntloadh , \SAEXE/RFIO/phrefendh , \SAEXE/RFIO/RIN1TRS , 
        \SAEXE/RFIO/n380 , \SAEXE/RFIO/n401 , \SAEXE/RFIO/nfst[0] , 
        \SAEXE/RFIO/n359 , \SAEXE/RFIO/n365 , \SAEXE/RFIO/phrfin1sah , 
        \SAEXE/RFIO/rfin2h , \SAEXE/RFIO/n358 , \SAEXE/RFIO/n376 , 
        \SAEXE/RFIO/n393 , \SAEXE/RFIO/n388 , \SAEXE/RFIO/n381 , 
        \SAEXE/RFIO/n364 , \SAEXE/RFIO/fst[1] , \SAEXE/RFIO/n400 , 
        \SAEXE/RFIO/srcadr1_h , \SAEXE/RFIO/n386 , \SAEXE/RFIO/n407 , 
        \SAEXE/RFIO/n363 , \SAEXE/RFIO/n378 , \SAEXE/RFIO/fst[2] , 
        \SAEXE/RFIO/n354 , \SAEXE/RFIO/n356 , \SAEXE/RFIO/n371 , 
        \SAEXE/RFIO/n361 , \SAEXE/RFIO/n394 , \SAEXE/RFIO/n384 , 
        \SAEXE/RFIO/n405 , \SAEXE/RFIO/n396 , \SAEXE/RFIO/n373 , 
        \SAEXE/RFIO/n353 , \SAEXE/RFIO/n368 , \SAEXE/RFIO/n374 , 
        \SAEXE/RFIO/fst[0] , \SAEXE/RFIO/n391 , \SAEXE/RFIO/cnt4dech , 
        \SAEXE/RFIO/rfin1tpenh , \SAEXE/RFIO/phrfin1h , \SAEXE/RFIO/n383 , 
        \SAEXE/RFIO/n366 , \SAEXE/RFIO/n402 , \SAEXE/RFIO/n398 , 
        \SAEXE/RFIO/n375 , \SAEXE/RFIO/n390 , \SAEXE/RFIO/n352 , 
        \SAEXE/RFIO/nfst[1] , \SAEXE/RFIO/*cell*3735/U61/Z_0 , 
        \SAEXE/RFIO/n399 , \SAEXE/RFIO/n367 , \SAEXE/RFIO/cnt4out[1] , 
        \SAEXE/RFIO/n382 , \SAEXE/RFIO/n403 , \SAEXE/RFIO/n385 , 
        \SAEXE/RFIO/n404 , \SAEXE/RFIO/ri1_trscdech , \SAEXE/RFIO/n360 , 
        \SAEXE/RFIO/nfst[3] , \SAEXE/RFIO/rfio1h , \SAEXE/RFIO/n355 , 
        \SAEXE/RFIO/n369 , \SAEXE/RFIO/n372 , \SAEXE/RFIO/n397 , 
        \SADR/SELOPR/n10656 , \SADR/SELOPR/n10683 , \SADR/SELOPR/n10698 , 
        \SADR/SELOPR/n10708 , \SADR/SELOPR/n10713 , \SADR/SELOPR/n10666 , 
        \SADR/SELOPR/n10674 , \SADR/SELOPR/n10691 , \SADR/SELOPR/n10701 , 
        \SADR/SELOPR/n10726 , \SADR/SELOPR/n10668 , \SADR/SELOPR/n10673 , 
        \SADR/SELOPR/n10696 , \SADR/SELOPR/n10706 , \SADR/SELOPR/n10721 , 
        \SADR/SELOPR/n10661 , \SADR/SELOPR/n10672 , \SADR/SELOPR/n10684 , 
        \SADR/SELOPR/n10714 , \SADR/SELOPR/n10728 , \SADR/SELOPR/n10697 , 
        \SADR/SELOPR/n10707 , \SADR/SELOPR/n10720 , \SADR/SELOPR/n10669 , 
        \SADR/SELOPR/n10685 , \SADR/SELOPR/n10729 , \SADR/SELOPR/n10715 , 
        \SADR/SELOPR/n10660 , \SADR/SELOPR/n10667 , \SADR/SELOPR/n10682 , 
        \SADR/SELOPR/n10712 , \SADR/SELOPR/n10699 , \SADR/SELOPR/n10709 , 
        \SADR/SELOPR/n10659 , \SADR/SELOPR/n10675 , \SADR/SELOPR/n10690 , 
        \SADR/SELOPR/n10727 , \SADR/SELOPR/n10700 , \SADR/SELOPR/n10680 , 
        \SADR/SELOPR/n10710 , \SADR/SELOPR/n10665 , \SADR/SELOPR/n10677 , 
        \SADR/SELOPR/n10670 , \SADR/SELOPR/n10689 , \SADR/SELOPR/n10692 , 
        \SADR/SELOPR/n10702 , \SADR/SELOPR/n10725 , \SADR/SELOPR/n10695 , 
        \SADR/SELOPR/n10705 , \SADR/SELOPR/n10719 , \SADR/SELOPR/n10722 , 
        \SADR/SELOPR/n10657 , \SADR/SELOPR/n10662 , \SADR/SELOPR/n10730 , 
        \SADR/SELOPR/n10687 , \SADR/SELOPR/n10717 , \SADR/SELOPR/n10679 , 
        \SADR/SELOPR/n10671 , \SADR/SELOPR/n10678 , \SADR/SELOPR/n10694 , 
        \SADR/SELOPR/n10723 , \SADR/SELOPR/n10704 , \SADR/SELOPR/n10663 , 
        \SADR/SELOPR/n10686 , \SADR/SELOPR/n10716 , \SADR/SELOPR/n10664 , 
        \SADR/SELOPR/n10681 , \SADR/SELOPR/n10711 , \SADR/SELOPR/n10658 , 
        \SADR/SELOPR/n10688 , \SADR/SELOPR/n10718 , \SADR/SELOPR/n10693 , 
        \SADR/SELOPR/n10703 , \SADR/SELOPR/n10724 , \SADR/SELOPR/n10676 , 
        \SADR/MAINSADR/n8879 , \SADR/MAINSADR/oddadd[20] , 
        \SADR/MAINSADR/oddadd[13] , \SADR/MAINSADR/addindoff[23] , 
        \SADR/MAINSADR/addindoff[19] , \SADR/MAINSADR/addindoff[8] , 
        \SADR/MAINSADR/n8669 , \SADR/MAINSADR/n8797 , 
        \SADR/MAINSADR/oddadd_m1[14] , \SADR/MAINSADR/oddadd_p2[15] , 
        \SADR/MAINSADR/n8772 , \SADR/MAINSADR/n8830 , \SADR/MAINSADR/n8755 , 
        \SADR/MAINSADR/n8817 , \SADR/MAINSADR/addindoff[10] , 
        \SADR/MAINSADR/addindoff[1] , \SADR/MAINSADR/n8655 , 
        \SADR/MAINSADR/n8769 , \SADR/MAINSADR/n8917 , \SADR/MAINSADR/n8672 , 
        \SADR/MAINSADR/n8887 , \SADR/MAINSADR/n8697 , \SADR/MAINSADR/n8845 , 
        \SADR/MAINSADR/n8707 , \SADR/MAINSADR/n8720 , 
        \SADR/MAINSADR/oddadd_m1[23] , \SADR/MAINSADR/oddadd_m1[10] , 
        \SADR/MAINSADR/oddadd_p2[22] , \SADR/MAINSADR/n8857 , 
        \SADR/MAINSADR/n8862 , \SADR/MAINSADR/oddadd_p2[11] , 
        \SADR/MAINSADR/n8685 , \SADR/MAINSADR/n8715 , \SADR/MAINSADR/n8732 , 
        \SADR/MAINSADR/n8870 , \SADR/MAINSADR/n8647 , 
        \SADR/MAINSADR/oddadd[17] , \SADR/MAINSADR/n8895 , 
        \SADR/MAINSADR/n8905 , \SADR/MAINSADR/n8922 , \SADR/MAINSADR/n8747 , 
        \SADR/MAINSADR/n8660 , \SADR/MAINSADR/n8760 , \SADR/MAINSADR/n8839 , 
        \SADR/MAINSADR/n8805 , \SADR/MAINSADR/n8822 , 
        \SADR/MAINSADR/addindoff[16] , \SADR/MAINSADR/addindoff[14] , 
        \SADR/MAINSADR/oddadd_p2[18] , \SADR/MAINSADR/addindoff[5] , 
        \SADR/MAINSADR/n8785 , \SADR/MAINSADR/oddadd_m1[19] , 
        \SADR/MAINSADR/n8729 , \SADR/MAINSADR/n8635 , \SADR/MAINSADR/n8782 , 
        \SADR/MAINSADR/addindoff[7] , \SADR/MAINSADR/n8802 , 
        \SADR/MAINSADR/n8699 , \SADR/MAINSADR/n8709 , \SADR/MAINSADR/n8740 , 
        \SADR/MAINSADR/n8825 , \SADR/MAINSADR/n8767 , \SADR/MAINSADR/n8889 , 
        \SADR/MAINSADR/n8919 , \SADR/MAINSADR/addindoff[21] , 
        \SADR/MAINSADR/addindoff[12] , \SADR/MAINSADR/addindoff[3] , 
        \SADR/MAINSADR/oddadd[18] , \SADR/MAINSADR/oddadd[15] , 
        \SADR/MAINSADR/n8667 , \SADR/MAINSADR/n8640 , \SADR/MAINSADR/n8892 , 
        \SADR/MAINSADR/n8902 , \SADR/MAINSADR/n8925 , 
        \SADR/MAINSADR/oddadd_m1[21] , \SADR/MAINSADR/oddadd_m1[12] , 
        \SADR/MAINSADR/oddadd_p2[20] , \SADR/MAINSADR/n8819 , 
        \SADR/MAINSADR/n8877 , \SADR/MAINSADR/oddadd_p2[13] , 
        \SADR/MAINSADR/n8735 , \SADR/MAINSADR/n8682 , \SADR/MAINSADR/n8712 , 
        \SADR/MAINSADR/n8850 , \SADR/MAINSADR/n8799 , \SADR/MAINSADR/n8727 , 
        \SADR/MAINSADR/n8865 , \SADR/MAINSADR/n8690 , \SADR/MAINSADR/n8700 , 
        \SADR/MAINSADR/n8842 , \SADR/MAINSADR/n8749 , \SADR/MAINSADR/n8675 , 
        \SADR/MAINSADR/oddadd_m1[16] , \SADR/MAINSADR/n8649 , 
        \SADR/MAINSADR/n8652 , \SADR/MAINSADR/n8880 , \SADR/MAINSADR/n8910 , 
        \SADR/MAINSADR/n8752 , \SADR/MAINSADR/oddadd[22] , 
        \SADR/MAINSADR/oddadd_p2[17] , \SADR/MAINSADR/n8810 , 
        \SADR/MAINSADR/n8837 , \SADR/MAINSADR/n8775 , \SADR/MAINSADR/n8859 , 
        \SADR/MAINSADR/oddadd[11] , \SADR/MAINSADR/n8790 , 
        \SADR/MAINSADR/index[6] , \SADR/MAINSADR/n8734 , \SADR/MAINSADR/n8876 , 
        \SADR/MAINSADR/oddadd_p2[8] , \SADR/MAINSADR/n8683 , 
        \SADR/MAINSADR/n8713 , \SADR/MAINSADR/n8851 , 
        \SADR/MAINSADR/offset[14] , \SADR/MAINSADR/n8666 , 
        \SADR/MAINSADR/n8798 , \SADR/MAINSADR/n8924 , \SADR/MAINSADR/n8893 , 
        \SADR/MAINSADR/n8903 , \SADR/MAINSADR/n8641 , 
        \SADR/MAINSADR/offset[2] , \SADR/MAINSADR/index[15] , 
        \SADR/MAINSADR/oddadd_m1[4] , \SADR/MAINSADR/oddadd_m2[7] , 
        \SADR/MAINSADR/n8818 , \SADR/MAINSADR/oddadd_p1[21] , 
        \SADR/MAINSADR/oddadd_p1[12] , \SADR/MAINSADR/oddadd_p1[2] , 
        \SADR/MAINSADR/oddadd[3] , \SADR/MAINSADR/n8741 , 
        \SADR/MAINSADR/n8803 , \SADR/MAINSADR/n8824 , \SADR/MAINSADR/n8766 , 
        \SADR/MAINSADR/n8918 , \SADR/MAINSADR/n8888 , 
        \SADR/MAINSADR/oddadd_p2[1] , \SADR/MAINSADR/n8634 , 
        \SADR/MAINSADR/n8783 , \SADR/MAINSADR/oddadd_m2[20] , 
        \SADR/MAINSADR/oddadd_m2[13] , \SADR/MAINSADR/n8698 , 
        \SADR/MAINSADR/n8708 , \SADR/MAINSADR/index[22] , 
        \SADR/MAINSADR/index[11] , \SADR/MAINSADR/oddadd[7] , 
        \SADR/MAINSADR/n8858 , \SADR/MAINSADR/offset[6] , 
        \SADR/MAINSADR/oddadd_m1[0] , \SADR/MAINSADR/oddadd_m2[3] , 
        \SADR/MAINSADR/offset[23] , \SADR/MAINSADR/n8791 , 
        \SADR/MAINSADR/offset[10] , \SADR/MAINSADR/n8648 , 
        \SADR/MAINSADR/index[2] , \SADR/MAINSADR/n8753 , \SADR/MAINSADR/n8774 , 
        \SADR/MAINSADR/n8811 , \SADR/MAINSADR/n8836 , 
        \SADR/MAINSADR/index[18] , \SADR/MAINSADR/oddadd_p1[16] , 
        \SADR/MAINSADR/oddadd_p2[5] , \SADR/MAINSADR/oddadd_m2[17] , 
        \SADR/MAINSADR/n8748 , \SADR/MAINSADR/n8674 , \SADR/MAINSADR/n8881 , 
        \SADR/MAINSADR/n8911 , \SADR/MAINSADR/oddadd_p1[6] , 
        \SADR/MAINSADR/oddadd_m1[9] , \SADR/MAINSADR/n8653 , 
        \SADR/MAINSADR/offset[19] , \SADR/MAINSADR/n8691 , 
        \SADR/MAINSADR/n8864 , \SADR/MAINSADR/n8726 , \SADR/MAINSADR/n8701 , 
        \SADR/MAINSADR/oddadd_m2[8] , \SADR/MAINSADR/n8843 , 
        \SADR/MAINSADR/n8844 , \SADR/MAINSADR/n8696 , \SADR/MAINSADR/n8706 , 
        \SADR/MAINSADR/n8721 , \SADR/MAINSADR/n8863 , \SADR/MAINSADR/index[9] , 
        \SADR/MAINSADR/oddadd_p1[14] , \SADR/MAINSADR/oddadd_p1[4] , 
        \SADR/MAINSADR/oddadd_m2[15] , \SADR/MAINSADR/n8768 , 
        \SADR/MAINSADR/n8654 , \SADR/MAINSADR/n8886 , \SADR/MAINSADR/n8916 , 
        \SADR/MAINSADR/oddadd_p2[7] , \SADR/MAINSADR/n8668 , 
        \SADR/MAINSADR/n8673 , \SADR/MAINSADR/index[0] , 
        \SADR/MAINSADR/index[20] , \SADR/MAINSADR/n8754 , 
        \SADR/MAINSADR/n8773 , \SADR/MAINSADR/n8816 , \SADR/MAINSADR/n8831 , 
        \SADR/MAINSADR/n8878 , \SADR/MAINSADR/index[13] , 
        \SADR/MAINSADR/offset[4] , \SADR/MAINSADR/oddadd[5] , 
        \SADR/MAINSADR/oddadd_m2[1] , \SADR/MAINSADR/offset[21] , 
        \SADR/MAINSADR/oddadd_m1[2] , \SADR/MAINSADR/n8796 , 
        \SADR/MAINSADR/offset[12] , \SADR/MAINSADR/oddadd_p1[23] , 
        \SADR/MAINSADR/oddadd_p1[10] , \SADR/MAINSADR/oddadd_p2[3] , 
        \SADR/MAINSADR/oddadd_p1[0] , \SADR/MAINSADR/n8633 , 
        \SADR/MAINSADR/oddadd_m2[22] , \SADR/MAINSADR/n8784 , 
        \SADR/MAINSADR/oddadd[8] , \SADR/MAINSADR/oddadd_m2[11] , 
        \SADR/MAINSADR/n8728 , \SADR/MAINSADR/n8761 , \SADR/MAINSADR/n8823 , 
        \SADR/MAINSADR/n8804 , \SADR/MAINSADR/n8746 , 
        \SADR/MAINSADR/offset[16] , \SADR/MAINSADR/offset[9] , 
        \SADR/MAINSADR/n8646 , \SADR/MAINSADR/offset[0] , 
        \SADR/MAINSADR/n8894 , \SADR/MAINSADR/n8904 , \SADR/MAINSADR/n8923 , 
        \SADR/MAINSADR/n8661 , \SADR/MAINSADR/oddadd_m1[6] , 
        \SADR/MAINSADR/index[17] , \SADR/MAINSADR/oddadd_m2[5] , 
        \SADR/MAINSADR/oddadd[1] , \SADR/MAINSADR/n8838 , 
        \SADR/MAINSADR/index[4] , \SADR/MAINSADR/n8684 , \SADR/MAINSADR/n8856 , 
        \SADR/MAINSADR/n8714 , \SADR/MAINSADR/n8733 , 
        \SADR/MAINSADR/oddadd_p1[19] , \SADR/MAINSADR/n8871 , 
        \SADR/MAINSADR/oddadd_p1[9] , \SADR/MAINSADR/oddadd_m2[18] , 
        \SADR/MAINSADR/oddadd_p1[22] , \SADR/MAINSADR/oddadd_p1[11] , 
        \SADR/MAINSADR/n8794 , \SADR/MAINSADR/oddadd_p1[1] , 
        \SADR/MAINSADR/oddadd_p2[2] , \SADR/MAINSADR/oddadd_m2[10] , 
        \SADR/MAINSADR/n8738 , \SADR/MAINSADR/n8771 , \SADR/MAINSADR/n8756 , 
        \SADR/MAINSADR/n8814 , \SADR/MAINSADR/n8833 , 
        \SADR/MAINSADR/index[16] , \SADR/MAINSADR/offset[17] , 
        \SADR/MAINSADR/offset[8] , \SADR/MAINSADR/oddadd[9] , 
        \SADR/MAINSADR/n8671 , \SADR/MAINSADR/n8928 , \SADR/MAINSADR/n8656 , 
        \SADR/MAINSADR/n8884 , \SADR/MAINSADR/n8914 , \SADR/MAINSADR/n8828 , 
        \SADR/MAINSADR/oddadd[0] , \SADR/MAINSADR/oddadd_m2[4] , 
        \SADR/MAINSADR/offset[1] , \SADR/MAINSADR/index[5] , 
        \SADR/MAINSADR/oddadd_m1[7] , \SADR/MAINSADR/oddadd_p1[18] , 
        \SADR/MAINSADR/n8723 , \SADR/MAINSADR/oddadd_p1[8] , 
        \SADR/MAINSADR/oddadd_m2[19] , \SADR/MAINSADR/n8694 , 
        \SADR/MAINSADR/n8704 , \SADR/MAINSADR/n8846 , \SADR/MAINSADR/n8861 , 
        \SADR/MAINSADR/n8638 , \SADR/MAINSADR/oddadd_m2[9] , 
        \SADR/MAINSADR/n8731 , \SADR/MAINSADR/n8873 , \SADR/MAINSADR/n8854 , 
        \SADR/MAINSADR/n8686 , \SADR/MAINSADR/n8716 , \SADR/MAINSADR/index[8] , 
        \SADR/MAINSADR/oddadd_p1[15] , \SADR/MAINSADR/oddadd_p1[5] , 
        \SADR/MAINSADR/cmpflg , \SADR/MAINSADR/oddadd_m2[14] , 
        \SADR/MAINSADR/n8778 , \SADR/MAINSADR/oddadd_p2[6] , 
        \SADR/MAINSADR/n8921 , \SADR/MAINSADR/n8663 , \SADR/MAINSADR/n8644 , 
        \SADR/MAINSADR/n8896 , \SADR/MAINSADR/n8906 , \SADR/MAINSADR/index[1] , 
        \SADR/MAINSADR/n8678 , \SADR/MAINSADR/n8744 , \SADR/MAINSADR/n8806 , 
        \SADR/MAINSADR/n8763 , \SADR/MAINSADR/offset[5] , 
        \SADR/MAINSADR/n8821 , \SADR/MAINSADR/oddadd_m1[3] , 
        \SADR/MAINSADR/index[21] , \SADR/MAINSADR/oddadd_m2[0] , 
        \SADR/MAINSADR/index[12] , \SADR/MAINSADR/oddadd[4] , 
        \SADR/MAINSADR/n8868 , \SADR/MAINSADR/offset[20] , 
        \SADR/MAINSADR/offset[13] , \SADR/MAINSADR/n8786 , 
        \SADR/MAINSADR/offset[7] , \SADR/MAINSADR/index[23] , 
        \SADR/MAINSADR/oddadd_m1[1] , \SADR/MAINSADR/oddadd_m2[2] , 
        \SADR/MAINSADR/n8848 , \SADR/MAINSADR/index[10] , 
        \SADR/MAINSADR/offset[22] , \SADR/MAINSADR/oddadd[6] , 
        \SADR/MAINSADR/n8636 , \SADR/MAINSADR/offset[11] , 
        \SADR/MAINSADR/n8781 , \SADR/MAINSADR/oddadd_p1[7] , 
        \SADR/MAINSADR/n8743 , \SADR/MAINSADR/index[3] , \SADR/MAINSADR/n8658 , 
        \SADR/MAINSADR/n8764 , \SADR/MAINSADR/n8826 , \SADR/MAINSADR/n8801 , 
        \SADR/MAINSADR/oddadd_p1[17] , \SADR/MAINSADR/oddadd_m2[16] , 
        \SADR/MAINSADR/n8758 , \SADR/MAINSADR/index[19] , 
        \SADR/MAINSADR/oddadd_p2[4] , \SADR/MAINSADR/n8643 , 
        \SADR/MAINSADR/n8891 , \SADR/MAINSADR/n8901 , \SADR/MAINSADR/n8664 , 
        \SADR/MAINSADR/n8926 , \SADR/MAINSADR/index[7] , 
        \SADR/MAINSADR/offset[18] , \SADR/MAINSADR/oddadd_m1[8] , 
        \SADR/MAINSADR/n8711 , \SADR/MAINSADR/n8681 , \SADR/MAINSADR/n8853 , 
        \SADR/MAINSADR/n8874 , \SADR/MAINSADR/n8736 , \SADR/MAINSADR/n8693 , 
        \SADR/MAINSADR/n8703 , \SADR/MAINSADR/oddadd_p2[9] , 
        \SADR/MAINSADR/n8841 , \SADR/MAINSADR/n8724 , \SADR/MAINSADR/n8866 , 
        \SADR/MAINSADR/n8788 , \SADR/MAINSADR/index[14] , 
        \SADR/MAINSADR/offset[15] , \SADR/MAINSADR/n8651 , 
        \SADR/MAINSADR/n8883 , \SADR/MAINSADR/n8913 , \SADR/MAINSADR/n8676 , 
        \SADR/MAINSADR/oddadd[2] , \SADR/MAINSADR/n8808 , 
        \SADR/MAINSADR/offset[3] , \SADR/MAINSADR/oddadd_m2[6] , 
        \SADR/MAINSADR/oddadd_m1[5] , \SADR/MAINSADR/oddadd_p1[20] , 
        \SADR/MAINSADR/oddadd_p1[13] , \SADR/MAINSADR/oddadd_p1[3] , 
        \SADR/MAINSADR/n8834 , \SADR/MAINSADR/n8751 , \SADR/MAINSADR/n8776 , 
        \SADR/MAINSADR/n8813 , \SADR/MAINSADR/n8898 , \SADR/MAINSADR/n8908 , 
        \SADR/MAINSADR/oddadd_p2[0] , \SADR/MAINSADR/n8793 , 
        \SADR/MAINSADR/addindoff[20] , \SADR/MAINSADR/addindoff[13] , 
        \SADR/MAINSADR/addindoff[2] , \SADR/MAINSADR/oddadd[19] , 
        \SADR/MAINSADR/oddadd_m2[21] , \SADR/MAINSADR/oddadd_m2[12] , 
        \SADR/MAINSADR/n8688 , \SADR/MAINSADR/n8718 , \SADR/MAINSADR/n8680 , 
        \SADR/MAINSADR/n8710 , \SADR/MAINSADR/n8737 , \SADR/MAINSADR/n8852 , 
        \SADR/MAINSADR/n8875 , \SADR/MAINSADR/ovf_addindoff , 
        \SADR/MAINSADR/n8759 , \SADR/MAINSADR/n8642 , \SADR/MAINSADR/n8890 , 
        \SADR/MAINSADR/n8900 , \SADR/MAINSADR/n8665 , 
        \SADR/MAINSADR/oddadd_m1[17] , \SADR/MAINSADR/n8927 , 
        \SADR/MAINSADR/oddadd_p2[16] , \SADR/MAINSADR/n8659 , 
        \SADR/MAINSADR/n8827 , \SADR/MAINSADR/n8765 , \SADR/MAINSADR/n8742 , 
        \SADR/MAINSADR/n8800 , \SADR/MAINSADR/n8849 , 
        \SADR/MAINSADR/addindoff[17] , \SADR/MAINSADR/oddadd[23] , 
        \SADR/MAINSADR/n8637 , \SADR/MAINSADR/oddadd[10] , 
        \SADR/MAINSADR/n8780 , \SADR/MAINSADR/addindoff[6] , 
        \SADR/MAINSADR/n8792 , \SADR/MAINSADR/oddadd[14] , 
        \SADR/MAINSADR/n8750 , \SADR/MAINSADR/n8689 , \SADR/MAINSADR/n8719 , 
        \SADR/MAINSADR/n8777 , \SADR/MAINSADR/n8835 , \SADR/MAINSADR/n8812 , 
        \SADR/MAINSADR/n8650 , \SADR/MAINSADR/n8882 , \SADR/MAINSADR/n8899 , 
        \SADR/MAINSADR/n8909 , \SADR/MAINSADR/n8912 , \SADR/MAINSADR/n8677 , 
        \SADR/MAINSADR/oddadd[16] , \SADR/MAINSADR/oddadd_m1[22] , 
        \SADR/MAINSADR/oddadd_m1[20] , \SADR/MAINSADR/oddadd_m1[13] , 
        \SADR/MAINSADR/oddadd_p2[21] , \SADR/MAINSADR/n8692 , 
        \SADR/MAINSADR/n8702 , \SADR/MAINSADR/n8809 , \SADR/MAINSADR/n8840 , 
        \SADR/MAINSADR/oddadd_p2[12] , \SADR/MAINSADR/n8725 , 
        \SADR/MAINSADR/n8867 , \SADR/MAINSADR/n8789 , 
        \SADR/MAINSADR/oddadd_m1[11] , \SADR/MAINSADR/oddadd_p2[10] , 
        \SADR/MAINSADR/n8722 , \SADR/MAINSADR/n8847 , \SADR/MAINSADR/n8860 , 
        \SADR/MAINSADR/n8639 , \SADR/MAINSADR/n8695 , \SADR/MAINSADR/n8705 , 
        \SADR/MAINSADR/n8670 , \SADR/MAINSADR/n8657 , \SADR/MAINSADR/n8829 , 
        \SADR/MAINSADR/n8885 , \SADR/MAINSADR/n8915 , \SADR/MAINSADR/n8815 , 
        \SADR/MAINSADR/addindoff[15] , \SADR/MAINSADR/n8757 , 
        \SADR/MAINSADR/n8770 , \SADR/MAINSADR/n8832 , 
        \SADR/MAINSADR/addindoff[4] , \SADR/MAINSADR/oddadd_m1[18] , 
        \SADR/MAINSADR/oddadd_p2[19] , \SADR/MAINSADR/n8795 , 
        \SADR/MAINSADR/n8787 , \SADR/MAINSADR/n8739 , \SADR/MAINSADR/n8869 , 
        \SADR/MAINSADR/oddadd_p2[14] , \SADR/MAINSADR/addindoff[18] , 
        \SADR/MAINSADR/addindoff[9] , \SADR/MAINSADR/oddadd[21] , 
        \SADR/MAINSADR/oddadd[12] , \SADR/MAINSADR/oddadd_m1[15] , 
        \SADR/MAINSADR/n8679 , \SADR/MAINSADR/n8745 , \SADR/MAINSADR/n8807 , 
        \SADR/MAINSADR/addindoff[0] , \SADR/MAINSADR/n8762 , 
        \SADR/MAINSADR/n8820 , \SADR/MAINSADR/n8779 , \SADR/MAINSADR/n8920 , 
        \SADR/MAINSADR/addindoff[22] , \SADR/MAINSADR/addindoff[11] , 
        \SADR/MAINSADR/n8662 , \SADR/MAINSADR/n8645 , \SADR/MAINSADR/n8897 , 
        \SADR/MAINSADR/n8907 , \SADR/MAINSADR/n8687 , \SADR/MAINSADR/n8717 , 
        \SADR/MAINSADR/n8730 , \SADR/MAINSADR/n8855 , \SADR/MAINSADR/n8872 , 
        \REGF/pbmemff21/RO_PPC19B114[9] , \REGF/pbmemff21/RO_PC19B72[6] , 
        \REGF/pbmemff21/RO_PPC19B114[0] , \REGF/pbmemff21/RO_PC19B72[2] , 
        \REGF/pbmemff21/n_853 , \REGF/pbmemff21/RO_PPC19B114[4] , 
        \REGF/pbmemff21/RO_PC19B72[9] , \REGF/pbmemff21/RO_PPC19B114[6] , 
        \REGF/pbmemff21/n6970 , \REGF/pbmemff21/RO_PC19B72[0] , 
        \REGF/pbmemff21/RO_PPC19B114[2] , \REGF/pbmemff21/RO_PC19B72[4] , 
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 , 
        \REGF/pbmemff21/RO_PPC19B114[13] , \REGF/pbmemff21/RO_PC19B72[14] , 
        \REGF/pbmemff21/RO_PC19BT[13] , \REGF/pbmemff21/RO_PC19BT[2] , 
        \REGF/pbmemff21/RO_PC19B72[10] , \REGF/pbmemff21/RO_PC19BT[17] , 
        \REGF/pbmemff21/RO_PC19BT[6] , \REGF/pbmemff21/RO_PC19BT[15] , 
        \REGF/pbmemff21/RO_PC19BT[4] , \REGF/pbmemff21/n6971 , 
        \REGF/pbmemff21/RO_PPC19B114[17] , \REGF/pbmemff21/RO_PC19B72[16] , 
        \REGF/pbmemff21/RO_PPC19B114[15] , \REGF/pbmemff21/RO_PC19B72[12] , 
        \REGF/pbmemff21/RO_PPC19B114[11] , \REGF/pbmemff21/RO_PC19BT[9] , 
        \REGF/pbmemff21/RO_PPC19B114[18] , \REGF/pbmemff21/RO_PC19BT[11] , 
        \REGF/pbmemff21/RO_PC19BT[0] , \REGF/pbmemff21/RO_PC19BT[18] , 
        \REGF/pbmemff21/RO_PC19BT[10] , \REGF/pbmemff21/RO_PC19BT[1] , 
        \REGF/pbmemff21/RO_PPC19B114[10] , \REGF/pbmemff21/RO_PC19B72[17] , 
        \REGF/pbmemff21/RO_PC19B72[13] , \REGF/pbmemff21/RO_PC19BT[8] , 
        \REGF/pbmemff21/RO_PC19BT[14] , \REGF/pbmemff21/RO_PC19BT[5] , 
        \REGF/pbmemff21/RO_PPC19B114[14] , \REGF/pbmemff21/RO_PC19B72[11] , 
        \REGF/pbmemff21/RO_PC19BT[16] , \REGF/pbmemff21/RO_PC19BT[7] , 
        \REGF/pbmemff21/RO_PC19B72[15] , \REGF/pbmemff21/RO_PPC19B114[16] , 
        \REGF/pbmemff21/RO_PC19B72[18] , \REGF/pbmemff21/RO_PC19BT[12] , 
        \REGF/pbmemff21/RO_PC19BT[3] , \REGF/pbmemff21/RO_PPC19B114[12] , 
        \REGF/pbmemff21/RO_PPC19B114[3] , \REGF/pbmemff21/RO_PC19B72[5] , 
        \REGF/pbmemff21/n6969 , \REGF/pbmemff21/RO_PC19B72[8] , 
        \REGF/pbmemff21/RO_PPC19B114[7] , \REGF/pbmemff21/RO_PC19B72[1] , 
        \REGF/pbmemff21/RO_PC19B72[3] , \REGF/pbmemff21/RO_PPC19B114[5] , 
        \REGF/pbmemff21/RO_PPC19B114[8] , \REGF/pbmemff21/RO_PC19B72[7] , 
        \REGF/pbmemff21/RO_PPC19B114[1] , \REG_2/ph8dec_1/n23 , 
        \REG_2/ph8dec_1/n22 , \SADR/ADDIDX/pgovfwxyzT , 
        \SADR/ADDIDX/pgovfwxyT , \SADR/ADDIDX/pgovfwyzT , 
        \SADR/ADDIDX/pgovfwxzT , \SADR/ADDIDX/pgovfxyzT , \SAEXE/SRC2/nqst[0] , 
        \SAEXE/SRC2/n185 , \SAEXE/SRC2/n190 , \SAEXE/SRC2/nqst[3] , 
        \SAEXE/SRC2/n205 , \SAEXE/SRC2/n217 , \SAEXE/SRC2/n222 , 
        \SAEXE/SRC2/eqst[4] , \SAEXE/SRC2/n199 , \SAEXE/SRC2/n219 , 
        \SAEXE/SRC2/n184 , \SAEXE/SRC2/eqst[2] , \SAEXE/SRC2/nqst[1] , 
        \SAEXE/SRC2/n202 , \SAEXE/SRC2/n210 , \SAEXE/SRC2/n197 , 
        \SAEXE/SRC2/n203 , \SAEXE/SRC2/n186 , \SAEXE/SRC2/n188 , 
        \SAEXE/SRC2/n191 , \SAEXE/SRC2/n196 , \SAEXE/SRC2/n218 , 
        \SAEXE/SRC2/n211 , \SAEXE/SRC2/n216 , \SAEXE/SRC2/n193 , 
        \SAEXE/SRC2/n198 , \SAEXE/SRC2/n204 , \SAEXE/SRC2/n214 , 
        \SAEXE/SRC2/n206 , \SAEXE/SRC2/n221 , \SAEXE/SRC2/n201 , 
        \SAEXE/SRC2/n213 , \SAEXE/SRC2/n187 , \SAEXE/SRC2/n194 , 
        \SAEXE/SRC2/n200 , \SAEXE/SRC2/n208 , \SAEXE/SRC2/n195 , 
        \SAEXE/SRC2/n209 , \SAEXE/SRC2/n189 , \SAEXE/SRC2/nqst[2] , 
        \SAEXE/SRC2/n212 , \SAEXE/SRC2/n215 , \SAEXE/SRC2/n192 , 
        \SAEXE/SRC2/n207 , \SAEXE/SRC2/eqst[1] , \SAEXE/SRC2/n220 , 
        \MCD/rd_wt_2/n4377 , \MCD/rd_wt_2/n4389 , \MCD/rd_wt_2/n4408 , 
        \MCD/rd_wt_2/n4392 , \MCD/rd_wt_2/n4413 , \MCD/rd_wt_2/n4379 , 
        \MCD/rd_wt_2/n4380 , \MCD/rd_wt_2/n4401 , \MCD/rd_wt_2/n4368 , 
        \MCD/rd_wt_2/n4370 , \MCD/rd_wt_2/n4387 , \MCD/rd_wt_2/n4406 , 
        \MCD/rd_wt_2/n4395 , \MCD/rd_wt_2/n4414 , \MCD/rd_wt_2/n4386 , 
        \MCD/rd_wt_2/ciff , \MCD/rd_wt_2/n4407 , \MCD/rd_wt_2/n4371 , 
        \MCD/rd_wt_2/n4378 , \MCD/rd_wt_2/n4394 , \MCD/rd_wt_2/n4415 , 
        \MCD/rd_wt_2/n4376 , \MCD/rd_wt_2/n4388 , \MCD/rd_wt_2/n4393 , 
        \MCD/rd_wt_2/n4412 , \MCD/rd_wt_2/n4409 , \MCD/rd_wt_2/n4374 , 
        \MCD/rd_wt_2/bacc , \MCD/rd_wt_2/n4381 , \MCD/rd_wt_2/n4391 , 
        \MCD/rd_wt_2/n4400 , \MCD/rd_wt_2/n4410 , \MCD/rd_wt_2/n4383 , 
        \MCD/rd_wt_2/n4384 , \MCD/rd_wt_2/n4398 , \MCD/rd_wt_2/n4402 , 
        \MCD/rd_wt_2/n4405 , \MCD/rd_wt_2/n4373 , \MCD/rd_wt_2/n4396 , 
        \MCD/rd_wt_2/n4417 , \MCD/rd_wt_2/n4369 , \MCD/rd_wt_2/n4385 , 
        \MCD/rd_wt_2/n4404 , \MCD/rd_wt_2/n4372 , \MCD/rd_wt_2/n4397 , 
        \MCD/rd_wt_2/n4416 , \MCD/rd_wt_2/n4367 , \MCD/rd_wt_2/n4375 , 
        \MCD/rd_wt_2/n4382 , \MCD/rd_wt_2/n4390 , \MCD/rd_wt_2/n4411 , 
        \MCD/rd_wt_2/n4399 , \MCD/rd_wt_2/n4403 , \REGF/pbmemff41/n7102 , 
        \REGF/pbmemff41/n7089 , \REGF/pbmemff41/n7092 , 
        \REGF/pbmemff41/RO_PSAS9B551[3] , 
        \REGF/pbmemff41/*cell*5493/U12/DATA2_0 , \REGF/pbmemff41/n_2861 , 
        \REGF/pbmemff41/*cell*5493/U2/DATA2_0 , \REGF/pbmemff41/n7087 , 
        \REGF/pbmemff41/*cell*5493/U59/Z_0 , \REGF/pbmemff41/n7095 , 
        \REGF/pbmemff41/RO_PSAS9B551[5] , 
        \REGF/pbmemff41/*cell*5493/U16/DATA2_0 , 
        \REGF/pbmemff41/*cell*5493/U6/DATA2_0 , \REGF/pbmemff41/RO_TRCOT[9] , 
        \REGF/pbmemff41/n7086 , \REGF/pbmemff41/RO_TRCOT[0] , 
        \REGF/pbmemff41/RO_TRCOT[14] , \REGF/pbmemff41/RO_TRCOT[23] , 
        \REGF/pbmemff41/RO_TRCOT[10] , \REGF/pbmemff41/n8037 , 
        \REGF/pbmemff41/n7094 , \REGF/pbmemff41/RO_TRCOT[19] , 
        \REGF/pbmemff41/RO_TRCOT[4] , \REGF/pbmemff41/RO_TRCOT[6] , 
        \REGF/pbmemff41/n7093 , \REGF/pbmemff41/n7103 , 
        \REGF/pbmemff41/*cell*5493/U10/DATA2_0 , \REGF/pbmemff41/n7088 , 
        \REGF/pbmemff41/RO_TRCOT[21] , \REGF/pbmemff41/RO_TRCOT[12] , 
        \REGF/pbmemff41/RO_TRCOT[2] , \REGF/pbmemff41/RO_TRCOT[16] , 
        \REGF/pbmemff41/*cell*5493/U14/DATA2_0 , 
        \REGF/pbmemff41/*cell*5493/U4/DATA2_0 , 
        \REGF/pbmemff41/*cell*5493/U79/Z_0 , \REGF/pbmemff41/RO_TRCOT[3] , 
        \REGF/pbmemff41/*cell*5493/U29/CONTROL1 , 
        \REGF/pbmemff41/*cell*5493/U20/DATA2_0 , \REGF/pbmemff41/RO_TRCOT[17] , 
        \REGF/pbmemff41/n7091 , \REGF/pbmemff41/n7101 , 
        \REGF/pbmemff41/*cell*5493/U63/Z_0 , \REGF/pbmemff41/RO_TRCOT[7] , 
        \REGF/pbmemff41/n_2859 , \REGF/pbmemff41/*cell*5493/U24/DATA2_0 , 
        \REGF/pbmemff41/*cell*5493/U77/Z_0 , \REGF/pbmemff41/n7083 , 
        \REGF/pbmemff41/n7098 , \REGF/pbmemff41/RO_TRCOT[20] , 
        \REGF/pbmemff41/RO_TRCOT[13] , \REGF/pbmemff41/RO_TRCOT[22] , 
        \REGF/pbmemff41/RO_TRCOT[11] , \REGF/pbmemff41/*cell*5493/U69/Z_0 , 
        \REGF/pbmemff41/n7084 , \REGF/pbmemff41/RO_TRCOT[18] , 
        \REGF/pbmemff41/RO_TRCOT[5] , \REGF/pbmemff41/*cell*5493/U73/Z_0 , 
        \REGF/pbmemff41/*cell*5493/U67/Z_0 , \REGF/pbmemff41/RO_TRCOT[8] , 
        \REGF/pbmemff41/RO_TRCOT[15] , \REGF/pbmemff41/RO_TRCOT[1] , 
        \REGF/pbmemff41/n7096 , \REGF/pbmemff41/*cell*5493/U27/CONTROL1 , 
        \REGF/pbmemff41/n8035 , \REGF/pbmemff41/n7085 , 
        \REGF/pbmemff41/RO_PSAS9B551[4] , \REGF/pbmemff41/*cell*5493/U75/Z_0 , 
        \REGF/pbmemff41/*cell*5493/U22/DATA2_0 , \REGF/pbmemff41/n8034 , 
        \REGF/pbmemff41/RO_PSAS9B551[0] , \REGF/pbmemff41/*cell*5493/U61/Z_0 , 
        \REGF/pbmemff41/n7097 , \REGF/pbmemff41/*cell*5493/U81/Z_0 , 
        \REGF/pbmemff41/*cell*5493/U65/Z_0 , \REGF/pbmemff41/n7090 , 
        \REGF/pbmemff41/n7100 , \REGF/pbmemff41/RO_PSAS9B551[2] , 
        \REGF/pbmemff41/n7099 , \REGF/pbmemff41/n7082 , 
        \REGF/pbmemff41/*cell*5493/U71/Z_0 , 
        \REGF/pbmemff41/*cell*5493/U129/CONTROL1 , 
        \REGF/pbmemff41/*cell*5493/U18/DATA2_0 , 
        \REGF/pbmemff41/*cell*5493/U8/DATA2_0 , \REGF/pbmemff61/n6505 , 
        \REGF/pbmemff61/RO_EXCO16B882[3] , \REGF/pbmemff61/RO_EXCO16B882[1] , 
        \REGF/pbmemff61/n6502 , \REGF/pbmemff61/n6503 , \REGF/pbmemff61/n6504 , 
        \REGF/pbmemff61/n_4044 , \REGF/pbmemff61/n6506 , 
        \REGF/pbmemff61/n6933 , \REGF/pbmemff61/n6501 , 
        \REGF/pbmemff61/RO_EXCO16B882[0] , \REGF/pbmemff61/n6500 , 
        \REGF/pbmemff61/RO_EXCO16B882[2] , \CONS/gte_124/n15 , 
        \CONS/gte_124/n55 , \CONS/gte_124/n32 , \CONS/gte_124/n29 , 
        \CONS/gte_124/n47 , \CONS/gte_124/n60 , \CONS/gte_124/n40 , 
        \CONS/gte_124/n16 , \CONS/gte_124/n27 , \CONS/gte_124/n35 , 
        \CONS/gte_124/n49 , \CONS/gte_124/n52 , \CONS/gte_124/n34 , 
        \CONS/gte_124/n26 , \CONS/gte_124/n41 , \CONS/gte_124/n53 , 
        \CONS/gte_124/n48 , \CONS/gte_124/n46 , \CONS/gte_124/n54 , 
        \CONS/gte_124/n61 , \CONS/gte_124/n28 , \CONS/gte_124/n33 , 
        \CONS/gte_124/n38 , \CONS/gte_124/n56 , \CONS/gte_124/n17 , 
        \CONS/gte_124/n18 , \CONS/gte_124/n24 , \CONS/gte_124/n31 , 
        \CONS/gte_124/n36 , \CONS/gte_124/n43 , \CONS/gte_124/n44 , 
        \CONS/gte_124/n58 , \CONS/gte_124/n37 , \CONS/gte_124/n51 , 
        \CONS/gte_124/n59 , \CONS/gte_124/n42 , \CONS/gte_124/n19 , 
        \CONS/gte_124/n50 , \CONS/gte_124/n25 , \CONS/gte_124/n39 , 
        \CONS/gte_124/n45 , \CONS/gte_124/n57 , \CONS/gte_124/n62 , 
        \CONS/gte_124/n30 , \CODEIF/CNT/wpfcen , \CODEIF/CNT/n3802 , 
        \CODEIF/CNT/n3775 , \CODEIF/CNT/n3790 , \CODEIF/CNT/n3810 , 
        \CODEIF/CNT/n3837 , \CODEIF/CNT/cst[2] , \CODEIF/CNT/n3767 , 
        \CODEIF/CNT/n3825 , \CODEIF/CNT/n3782 , \CODEIF/CNT/n3799 , 
        \CODEIF/CNT/cst[4] , \CODEIF/CNT/n3819 , \CODEIF/CNT/n3839 , 
        \CODEIF/CNT/n3805 , \CODEIF/CNT/n3785 , \CODEIF/CNT/n3822 , 
        \CODEIF/CNT/n3768 , \CODEIF/CNT/n3804 , \CODEIF/CNT/n3769 , 
        \CODEIF/CNT/n3772 , \CODEIF/CNT/n3797 , \CODEIF/CNT/n3817 , 
        \CODEIF/CNT/n3830 , \CODEIF/CNT/cst[0] , \CODEIF/CNT/n3823 , 
        \CODEIF/CNT/nst[3] , \CODEIF/CNT/n3784 , \CODEIF/CNT/n3838 , 
        \CODEIF/CNT/n3783 , \CODEIF/CNT/wwbregen , \CODEIF/CNT/n3773 , 
        \CODEIF/CNT/n3796 , \CODEIF/CNT/n3774 , \CODEIF/CNT/n3811 , 
        \CODEIF/CNT/n3816 , \CODEIF/CNT/n3831 , \CODEIF/CNT/n3836 , 
        \CODEIF/CNT/n3791 , \CODEIF/CNT/nst[1] , \CODEIF/CNT/n3798 , 
        \CODEIF/CNT/n3818 , \CODEIF/CNT/n3766 , \CODEIF/CNT/n3803 , 
        \CODEIF/CNT/n3824 , \CODEIF/CNT/n3808 , \CODEIF/CNT/n3806 , 
        \CODEIF/CNT/n3801 , \CODEIF/CNT/nst[0] , \CODEIF/CNT/n3788 , 
        \CODEIF/CNT/n3793 , \CODEIF/CNT/n3841 , \CODEIF/CNT/n3776 , 
        \CODEIF/CNT/n3834 , \CODEIF/CNT/n3813 , \CODEIF/CNT/n3826 , 
        \CODEIF/CNT/n3786 , \CODEIF/CNT/n3778 , \CODEIF/CNT/n3781 , 
        \CODEIF/CNT/nst[4] , \CODEIF/CNT/n3807 , \CODEIF/CNT/n3771 , 
        \CODEIF/CNT/n3814 , \CODEIF/CNT/n3821 , \CODEIF/CNT/nst[2] , 
        \CODEIF/CNT/n3794 , \CODEIF/CNT/n3833 , \CODEIF/CNT/n3828 , 
        \CODEIF/CNT/cst[1] , \CODEIF/CNT/n3820 , \CODEIF/CNT/n3779 , 
        \CODEIF/CNT/n3787 , \CODEIF/CNT/n3829 , \CODEIF/CNT/n3770 , 
        \CODEIF/CNT/n3795 , \CODEIF/CNT/n3815 , \CODEIF/CNT/n3777 , 
        \CODEIF/CNT/n3832 , \CODEIF/CNT/n3835 , \CODEIF/CNT/n3780 , 
        \CODEIF/CNT/n3789 , \CODEIF/CNT/n3792 , \CODEIF/CNT/n3812 , 
        \CODEIF/CNT/n3809 , \CODEIF/CNT/n3840 , \CODEIF/CNT/cst[3] , 
        \CODEIF/CNT/n3800 , \CODEIF/CNT/n3827 , \REGF/pbmemout1/n5695 , 
        \REGF/pbmemout1/n5705 , \REGF/pbmemout1/n5722 , \REGF/pbmemout1/n5860 , 
        \REGF/pbmemout1/n6233 , \REGF/pbmemout1/n6093 , \REGF/pbmemout1/n6103 , 
        \REGF/pbmemout1/n6124 , \REGF/pbmemout1/n5847 , \REGF/pbmemout1/n6214 , 
        \REGF/pbmemout1/n6384 , \REGF/pbmemout1/n6328 , \REGF/pbmemout1/n6018 , 
        \REGF/pbmemout1/n6188 , \REGF/pbmemout1/n5829 , \REGF/pbmemout1/n5932 , 
        \REGF/pbmemout1/n6051 , \REGF/pbmemout1/n5885 , \REGF/pbmemout1/n6361 , 
        \REGF/pbmemout1/n5915 , \REGF/pbmemout1/n6346 , \REGF/pbmemout1/n6076 , 
        \REGF/pbmemout1/n5757 , \REGF/pbmemout1/n5770 , \REGF/pbmemout1/n5815 , 
        \REGF/pbmemout1/n6176 , \REGF/pbmemout1/n5832 , \REGF/pbmemout1/n5985 , 
        \REGF/pbmemout1/n6246 , \REGF/pbmemout1/n6261 , \REGF/pbmemout1/n6151 , 
        \REGF/pbmemout1/n5739 , \REGF/pbmemout1/n5795 , \REGF/pbmemout1/n5929 , 
        \REGF/pbmemout1/n6284 , \REGF/pbmemout1/n6314 , \REGF/pbmemout1/n5947 , 
        \REGF/pbmemout1/n6024 , \REGF/pbmemout1/n6003 , \REGF/pbmemout1/n6193 , 
        \REGF/pbmemout1/n6333 , \REGF/pbmemout1/n5960 , \REGF/pbmemout1/n6088 , 
        \REGF/pbmemout1/n6118 , \REGF/pbmemout1/n6228 , \REGF/pbmemout1/n5787 , 
        \REGF/pbmemout1/n5869 , \REGF/pbmemout1/n6296 , \REGF/pbmemout1/n6306 , 
        \REGF/pbmemout1/n5955 , \REGF/pbmemout1/n6036 , \REGF/pbmemout1/n6181 , 
        \REGF/pbmemout1/n6011 , \REGF/pbmemout1/n5679 , \REGF/pbmemout1/n6321 , 
        \REGF/pbmemout1/n5972 , \REGF/pbmemout1/n6368 , \REGF/pbmemout1/n6058 , 
        \REGF/pbmemout1/n5745 , \REGF/pbmemout1/n5762 , \REGF/pbmemout1/n5807 , 
        \REGF/pbmemout1/n6164 , \REGF/pbmemout1/n5997 , \REGF/pbmemout1/n5820 , 
        \REGF/pbmemout1/n6254 , \REGF/pbmemout1/n6273 , \REGF/pbmemout1/n5779 , 
        \REGF/pbmemout1/n6143 , \REGF/pbmemout1/n6158 , \REGF/pbmemout1/n6268 , 
        \REGF/pbmemout1/n6043 , \REGF/pbmemout1/n5920 , \REGF/pbmemout1/n6373 , 
        \REGF/pbmemout1/n5897 , \REGF/pbmemout1/n5907 , \REGF/pbmemout1/n6354 , 
        \REGF/pbmemout1/n6064 , \REGF/pbmemout1/n5969 , \REGF/pbmemout1/n5687 , 
        \REGF/pbmemout1/n5730 , \REGF/pbmemout1/n5872 , \REGF/pbmemout1/n6221 , 
        \REGF/pbmemout1/n6111 , \REGF/pbmemout1/n6081 , \REGF/pbmemout1/n6136 , 
        \REGF/pbmemout1/n5717 , \REGF/pbmemout1/n5855 , \REGF/pbmemout1/n6206 , 
        \REGF/pbmemout1/n5949 , \REGF/pbmemout1/n5680 , \REGF/pbmemout1/n5710 , 
        \REGF/pbmemout1/n5852 , \REGF/pbmemout1/n6201 , \REGF/pbmemout1/n5737 , 
        \REGF/pbmemout1/n6131 , \REGF/pbmemout1/n5759 , \REGF/pbmemout1/n5875 , 
        \REGF/pbmemout1/n6086 , \REGF/pbmemout1/n6116 , \REGF/pbmemout1/n6226 , 
        \REGF/pbmemout1/n6178 , \REGF/pbmemout1/n6248 , \REGF/pbmemout1/n6063 , 
        \REGF/pbmemout1/n5742 , \REGF/pbmemout1/n5765 , \REGF/pbmemout1/n6353 , 
        \REGF/pbmemout1/n5890 , \REGF/pbmemout1/n5900 , \REGF/pbmemout1/n6374 , 
        \REGF/pbmemout1/n5927 , \REGF/pbmemout1/n6044 , \REGF/pbmemout1/n6348 , 
        \REGF/pbmemout1/n6078 , \REGF/pbmemout1/n6144 , \REGF/pbmemout1/n5800 , 
        \REGF/pbmemout1/n5827 , \REGF/pbmemout1/n6274 , \REGF/pbmemout1/n6253 , 
        \REGF/pbmemout1/n5990 , \REGF/pbmemout1/n6163 , \REGF/pbmemout1/n5849 , 
        \REGF/pbmemout1/n5975 , \REGF/pbmemout1/n6326 , \REGF/pbmemout1/n6016 , 
        \REGF/pbmemout1/n6186 , \REGF/pbmemout1/n5689 , \REGF/pbmemout1/n5780 , 
        \REGF/pbmemout1/n5792 , \REGF/pbmemout1/n5952 , \REGF/pbmemout1/n6031 , 
        \REGF/pbmemout1/n6291 , \REGF/pbmemout1/n6301 , \REGF/pbmemout1/n5967 , 
        \REGF/pbmemout1/n6334 , \REGF/pbmemout1/n6004 , \REGF/pbmemout1/n6194 , 
        \REGF/pbmemout1/n6023 , \REGF/pbmemout1/n5940 , \REGF/pbmemout1/n6283 , 
        \REGF/pbmemout1/n6313 , \REGF/pbmemout1/n6138 , \REGF/pbmemout1/n5719 , 
        \REGF/pbmemout1/n5750 , \REGF/pbmemout1/n5777 , \REGF/pbmemout1/n6208 , 
        \REGF/pbmemout1/n6156 , \REGF/pbmemout1/n5812 , \REGF/pbmemout1/n5835 , 
        \REGF/pbmemout1/n6266 , \REGF/pbmemout1/n6241 , \REGF/pbmemout1/n5982 , 
        \REGF/pbmemout1/n6171 , \REGF/pbmemout1/n5899 , \REGF/pbmemout1/n5909 , 
        \REGF/pbmemout1/n6071 , \REGF/pbmemout1/n5677 , \REGF/pbmemout1/n6341 , 
        \REGF/pbmemout1/n5882 , \REGF/pbmemout1/n5912 , \REGF/pbmemout1/n6366 , 
        \REGF/pbmemout1/n5935 , \REGF/pbmemout1/n6056 , \REGF/pbmemout1/n5809 , 
        \REGF/pbmemout1/n5999 , \REGF/pbmemout1/n5692 , \REGF/pbmemout1/n5840 , 
        \REGF/pbmemout1/n6213 , \REGF/pbmemout1/n6383 , \REGF/pbmemout1/n5702 , 
        \REGF/pbmemout1/n5725 , \REGF/pbmemout1/n6123 , \REGF/pbmemout1/n5789 , 
        \REGF/pbmemout1/n5867 , \REGF/pbmemout1/n6094 , \REGF/pbmemout1/n6104 , 
        \REGF/pbmemout1/n6234 , \REGF/pbmemout1/n6298 , \REGF/pbmemout1/n6308 , 
        \REGF/pbmemout1/n6038 , \REGF/pbmemout1/n5781 , \REGF/pbmemout1/n5848 , 
        \REGF/pbmemout1/n5974 , \REGF/pbmemout1/n6327 , \REGF/pbmemout1/n6017 , 
        \REGF/pbmemout1/n6187 , \REGF/pbmemout1/n6030 , \REGF/pbmemout1/n6290 , 
        \REGF/pbmemout1/n6300 , \REGF/pbmemout1/n5953 , \REGF/pbmemout1/n5743 , 
        \REGF/pbmemout1/O_LDO[27] , \REGF/pbmemout1/O_LDO[14] , 
        \REGF/pbmemout1/n6349 , \REGF/pbmemout1/n6079 , \REGF/pbmemout1/n5764 , 
        \REGF/pbmemout1/n5801 , \REGF/pbmemout1/n5826 , \REGF/pbmemout1/n6145 , 
        \REGF/pbmemout1/n6275 , \REGF/pbmemout1/n5991 , \REGF/pbmemout1/n6252 , 
        \REGF/pbmemout1/n5758 , \REGF/pbmemout1/n6162 , \REGF/pbmemout1/n6179 , 
        \REGF/pbmemout1/n6249 , \REGF/pbmemout1/O_LDO[7] , 
        \REGF/pbmemout1/n6062 , \REGF/pbmemout1/n5891 , \REGF/pbmemout1/n5901 , 
        \REGF/pbmemout1/n6352 , \REGF/pbmemout1/n5926 , \REGF/pbmemout1/n6375 , 
        \REGF/pbmemout1/n6045 , \REGF/pbmemout1/n5948 , \REGF/pbmemout1/n5681 , 
        \REGF/pbmemout1/n5853 , \REGF/pbmemout1/n6200 , \REGF/pbmemout1/n6130 , 
        \REGF/pbmemout1/n5703 , \REGF/pbmemout1/n5711 , \REGF/pbmemout1/n5736 , 
        \REGF/pbmemout1/n6087 , \REGF/pbmemout1/n6117 , \REGF/pbmemout1/n5841 , 
        \REGF/pbmemout1/n5874 , \REGF/pbmemout1/n6227 , \REGF/pbmemout1/n6212 , 
        \REGF/pbmemout1/n6382 , \REGF/pbmemout1/n6122 , \REGF/pbmemout1/n5693 , 
        \REGF/pbmemout1/n5724 , \REGF/pbmemout1/n6095 , \REGF/pbmemout1/n6105 , 
        \REGF/pbmemout1/O_LDO[23] , \REGF/pbmemout1/n5866 , 
        \REGF/pbmemout1/n6235 , \REGF/pbmemout1/n6299 , \REGF/pbmemout1/n6309 , 
        \REGF/pbmemout1/O_LDO[10] , \REGF/pbmemout1/n5788 , 
        \REGF/pbmemout1/n6039 , \REGF/pbmemout1/n6070 , \REGF/pbmemout1/n5883 , 
        \REGF/pbmemout1/n5913 , \REGF/pbmemout1/n6340 , \REGF/pbmemout1/n5934 , 
        \REGF/pbmemout1/n6367 , \REGF/pbmemout1/n6057 , \REGF/pbmemout1/n5808 , 
        \REGF/pbmemout1/n5998 , \REGF/pbmemout1/n5751 , \REGF/pbmemout1/n5776 , 
        \REGF/pbmemout1/n5813 , \REGF/pbmemout1/n5834 , \REGF/pbmemout1/n6157 , 
        \REGF/pbmemout1/n6267 , \REGF/pbmemout1/n5983 , \REGF/pbmemout1/n6240 , 
        \REGF/pbmemout1/n6170 , \REGF/pbmemout1/n5898 , \REGF/pbmemout1/n5908 , 
        \REGF/pbmemout1/O_LDO[3] , \REGF/pbmemout1/n6335 , 
        \REGF/pbmemout1/n5966 , \REGF/pbmemout1/n6005 , \REGF/pbmemout1/n6195 , 
        \REGF/pbmemout1/n5793 , \REGF/pbmemout1/n6022 , \REGF/pbmemout1/n6282 , 
        \REGF/pbmemout1/n6312 , \REGF/pbmemout1/n5941 , \REGF/pbmemout1/n5688 , 
        \REGF/pbmemout1/n5718 , \REGF/pbmemout1/O_LDO[19] , 
        \REGF/pbmemout1/n6139 , \REGF/pbmemout1/O_LDO[1] , 
        \REGF/pbmemout1/n5794 , \REGF/pbmemout1/n6209 , \REGF/pbmemout1/n5946 , 
        \REGF/pbmemout1/n6285 , \REGF/pbmemout1/n6315 , \REGF/pbmemout1/n6025 , 
        \REGF/pbmemout1/n6192 , \REGF/pbmemout1/n6002 , \REGF/pbmemout1/n5961 , 
        \REGF/pbmemout1/n6332 , \REGF/pbmemout1/n5738 , \REGF/pbmemout1/n6089 , 
        \REGF/pbmemout1/n6119 , \REGF/pbmemout1/O_LDO[31] , 
        \REGF/pbmemout1/n6229 , \REGF/pbmemout1/O_LDO[28] , 
        \REGF/pbmemout1/n5756 , \REGF/pbmemout1/n6177 , \REGF/pbmemout1/n5771 , 
        \REGF/pbmemout1/n5814 , \REGF/pbmemout1/n5984 , \REGF/pbmemout1/n6247 , 
        \REGF/pbmemout1/n5833 , \REGF/pbmemout1/n6260 , \REGF/pbmemout1/n6150 , 
        \REGF/pbmemout1/n5928 , \REGF/pbmemout1/n6050 , \REGF/pbmemout1/n6360 , 
        \REGF/pbmemout1/n5884 , \REGF/pbmemout1/n5914 , \REGF/pbmemout1/n5933 , 
        \REGF/pbmemout1/n6347 , \REGF/pbmemout1/n6077 , \REGF/pbmemout1/n5828 , 
        \REGF/pbmemout1/n5723 , \REGF/pbmemout1/n5861 , \REGF/pbmemout1/n6232 , 
        \REGF/pbmemout1/n5694 , \REGF/pbmemout1/n6102 , \REGF/pbmemout1/n6092 , 
        \REGF/pbmemout1/n5704 , \REGF/pbmemout1/O_LDO[21] , 
        \REGF/pbmemout1/O_LDO[8] , \REGF/pbmemout1/n5846 , 
        \REGF/pbmemout1/n6125 , \REGF/pbmemout1/n6215 , 
        \REGF/pbmemout1/O_LDO[12] , \REGF/pbmemout1/n6329 , 
        \REGF/pbmemout1/n6019 , \REGF/pbmemout1/n6189 , \REGF/pbmemout1/n5968 , 
        \REGF/pbmemout1/n5686 , \REGF/pbmemout1/n5716 , \REGF/pbmemout1/n5731 , 
        \REGF/pbmemout1/n5873 , \REGF/pbmemout1/n6220 , \REGF/pbmemout1/n6080 , 
        \REGF/pbmemout1/n6110 , \REGF/pbmemout1/O_LDO[5] , 
        \REGF/pbmemout1/n5778 , \REGF/pbmemout1/n5854 , \REGF/pbmemout1/n6137 , 
        \REGF/pbmemout1/n6207 , \REGF/pbmemout1/n6159 , \REGF/pbmemout1/n6269 , 
        \REGF/pbmemout1/n6042 , \REGF/pbmemout1/n6372 , \REGF/pbmemout1/n5921 , 
        \REGF/pbmemout1/n5896 , \REGF/pbmemout1/n6355 , \REGF/pbmemout1/n5906 , 
        \REGF/pbmemout1/n6065 , \REGF/pbmemout1/n5744 , \REGF/pbmemout1/n5678 , 
        \REGF/pbmemout1/O_LDO[25] , \REGF/pbmemout1/n6369 , 
        \REGF/pbmemout1/O_LDO[16] , \REGF/pbmemout1/n6059 , 
        \REGF/pbmemout1/n6165 , \REGF/pbmemout1/n5763 , \REGF/pbmemout1/n5806 , 
        \REGF/pbmemout1/n6255 , \REGF/pbmemout1/n5821 , \REGF/pbmemout1/n5996 , 
        \REGF/pbmemout1/n6272 , \REGF/pbmemout1/n6142 , \REGF/pbmemout1/n5786 , 
        \REGF/pbmemout1/n5868 , \REGF/pbmemout1/n5954 , \REGF/pbmemout1/n6297 , 
        \REGF/pbmemout1/n6307 , \REGF/pbmemout1/n6037 , \REGF/pbmemout1/n6010 , 
        \REGF/pbmemout1/n6180 , \REGF/pbmemout1/n5973 , \REGF/pbmemout1/n6320 , 
        \REGF/pbmemout1/n5978 , \REGF/pbmemout1/n5696 , \REGF/pbmemout1/n6127 , 
        \REGF/pbmemout1/n5706 , \REGF/pbmemout1/n5721 , \REGF/pbmemout1/n5844 , 
        \REGF/pbmemout1/n6217 , \REGF/pbmemout1/n5863 , \REGF/pbmemout1/n6230 , 
        \REGF/pbmemout1/n6100 , \REGF/pbmemout1/n6090 , 
        \REGF/pbmemout1/O_LDO[24] , \REGF/pbmemout1/O_LDO[4] , 
        \REGF/pbmemout1/n5768 , \REGF/pbmemout1/n6149 , \REGF/pbmemout1/n6279 , 
        \REGF/pbmemout1/n5916 , \REGF/pbmemout1/n5886 , \REGF/pbmemout1/n6345 , 
        \REGF/pbmemout1/n6075 , \REGF/pbmemout1/n6052 , \REGF/pbmemout1/n5931 , 
        \REGF/pbmemout1/n6362 , \REGF/pbmemout1/O_LDO[17] , 
        \REGF/pbmemout1/n6379 , \REGF/pbmemout1/n6049 , \REGF/pbmemout1/n5831 , 
        \REGF/pbmemout1/n6262 , \REGF/pbmemout1/n5754 , \REGF/pbmemout1/n5773 , 
        \REGF/pbmemout1/n6152 , \REGF/pbmemout1/n5816 , \REGF/pbmemout1/n6175 , 
        \REGF/pbmemout1/n5986 , \REGF/pbmemout1/n6245 , \REGF/pbmemout1/n5878 , 
        \REGF/pbmemout1/n5728 , \REGF/pbmemout1/O_LDO[0] , 
        \REGF/pbmemout1/n5796 , \REGF/pbmemout1/n6000 , \REGF/pbmemout1/n6190 , 
        \REGF/pbmemout1/n5963 , \REGF/pbmemout1/n6330 , \REGF/pbmemout1/n6287 , 
        \REGF/pbmemout1/n6317 , \REGF/pbmemout1/n5944 , \REGF/pbmemout1/n6027 , 
        \REGF/pbmemout1/n6012 , \REGF/pbmemout1/n6182 , \REGF/pbmemout1/n6322 , 
        \REGF/pbmemout1/n5971 , \REGF/pbmemout1/n6295 , \REGF/pbmemout1/n6305 , 
        \REGF/pbmemout1/n5956 , \REGF/pbmemout1/n5784 , \REGF/pbmemout1/n6035 , 
        \REGF/pbmemout1/O_LDO[30] , \REGF/pbmemout1/O_LDO[29] , 
        \REGF/pbmemout1/n6099 , \REGF/pbmemout1/n6109 , \REGF/pbmemout1/n6239 , 
        \REGF/pbmemout1/n5746 , \REGF/pbmemout1/n5761 , \REGF/pbmemout1/n5823 , 
        \REGF/pbmemout1/n6270 , \REGF/pbmemout1/n6140 , \REGF/pbmemout1/n5804 , 
        \REGF/pbmemout1/n6167 , \REGF/pbmemout1/n5994 , \REGF/pbmemout1/n6257 , 
        \REGF/pbmemout1/n5938 , \REGF/pbmemout1/n5894 , \REGF/pbmemout1/n5904 , 
        \REGF/pbmemout1/n6357 , \REGF/pbmemout1/n6067 , \REGF/pbmemout1/n6040 , 
        \REGF/pbmemout1/n5923 , \REGF/pbmemout1/n6370 , \REGF/pbmemout1/n5838 , 
        \REGF/pbmemout1/n5684 , \REGF/pbmemout1/n5714 , 
        \REGF/pbmemout1/O_LDO[9] , \REGF/pbmemout1/n6135 , 
        \REGF/pbmemout1/n5856 , \REGF/pbmemout1/n6205 , \REGF/pbmemout1/n5871 , 
        \REGF/pbmemout1/n6222 , \REGF/pbmemout1/n6082 , \REGF/pbmemout1/n6112 , 
        \REGF/pbmemout1/n5733 , \REGF/pbmemout1/n5683 , \REGF/pbmemout1/n5734 , 
        \REGF/pbmemout1/O_LDO[20] , \REGF/pbmemout1/n6339 , 
        \REGF/pbmemout1/O_LDO[13] , \REGF/pbmemout1/n6009 , 
        \REGF/pbmemout1/n6199 , \REGF/pbmemout1/n5851 , \REGF/pbmemout1/n5876 , 
        \REGF/pbmemout1/n6085 , \REGF/pbmemout1/n6115 , \REGF/pbmemout1/n6225 , 
        \REGF/pbmemout1/n6202 , \REGF/pbmemout1/n5713 , \REGF/pbmemout1/n6132 , 
        \REGF/pbmemout1/O_LDO[22] , \REGF/pbmemout1/O_LDO[11] , 
        \REGF/pbmemout1/n6289 , \REGF/pbmemout1/n6319 , \REGF/pbmemout1/n6029 , 
        \REGF/pbmemout1/n5798 , \REGF/pbmemout1/n6377 , \REGF/pbmemout1/n5924 , 
        \REGF/pbmemout1/n6047 , \REGF/pbmemout1/n6060 , \REGF/pbmemout1/n6350 , 
        \REGF/pbmemout1/n5893 , \REGF/pbmemout1/n5903 , \REGF/pbmemout1/n5741 , 
        \REGF/pbmemout1/n5803 , \REGF/pbmemout1/n5818 , \REGF/pbmemout1/n5988 , 
        \REGF/pbmemout1/n6250 , \REGF/pbmemout1/n5993 , \REGF/pbmemout1/n6160 , 
        \REGF/pbmemout1/n5766 , \REGF/pbmemout1/n6147 , \REGF/pbmemout1/n5824 , 
        \REGF/pbmemout1/n6277 , \REGF/pbmemout1/n5888 , \REGF/pbmemout1/n5918 , 
        \REGF/pbmemout1/n5698 , \REGF/pbmemout1/O_LDO[18] , 
        \REGF/pbmemout1/O_LDO[2] , \REGF/pbmemout1/n5783 , 
        \REGF/pbmemout1/n6032 , \REGF/pbmemout1/n5951 , \REGF/pbmemout1/n6302 , 
        \REGF/pbmemout1/n6292 , \REGF/pbmemout1/n5976 , \REGF/pbmemout1/n6325 , 
        \REGF/pbmemout1/n6015 , \REGF/pbmemout1/n6185 , \REGF/pbmemout1/n6129 , 
        \REGF/pbmemout1/n5708 , \REGF/pbmemout1/n6219 , \REGF/pbmemout1/n5858 , 
        \REGF/pbmemout1/O_LDO[26] , \REGF/pbmemout1/n5791 , 
        \REGF/pbmemout1/n6020 , \REGF/pbmemout1/n5943 , \REGF/pbmemout1/n6280 , 
        \REGF/pbmemout1/n6310 , \REGF/pbmemout1/n5964 , \REGF/pbmemout1/n6337 , 
        \REGF/pbmemout1/n6007 , \REGF/pbmemout1/n6197 , \REGF/pbmemout1/n6359 , 
        \REGF/pbmemout1/O_LDO[15] , \REGF/pbmemout1/n6069 , 
        \REGF/pbmemout1/n5811 , \REGF/pbmemout1/n6242 , \REGF/pbmemout1/n5981 , 
        \REGF/pbmemout1/n6172 , \REGF/pbmemout1/O_LDO[6] , 
        \REGF/pbmemout1/n5748 , \REGF/pbmemout1/n5753 , \REGF/pbmemout1/n5774 , 
        \REGF/pbmemout1/n6155 , \REGF/pbmemout1/n5836 , \REGF/pbmemout1/n6265 , 
        \REGF/pbmemout1/n6169 , \REGF/pbmemout1/n6259 , \REGF/pbmemout1/n6365 , 
        \REGF/pbmemout1/n5936 , \REGF/pbmemout1/n6055 , \REGF/pbmemout1/n6072 , 
        \REGF/pbmemout1/n6342 , \REGF/pbmemout1/n5881 , \REGF/pbmemout1/n5911 , 
        \REGF/pbmemout1/n5958 , \REGF/pbmemout1/n5691 , \REGF/pbmemout1/n5701 , 
        \REGF/pbmemout1/n5726 , \REGF/pbmemout1/n5843 , \REGF/pbmemout1/n5864 , 
        \REGF/pbmemout1/n6097 , \REGF/pbmemout1/n6107 , \REGF/pbmemout1/n6237 , 
        \REGF/pbmemout1/n6210 , \REGF/pbmemout1/n6380 , \REGF/pbmemout1/n5699 , 
        \REGF/pbmemout1/n5709 , \REGF/pbmemout1/n5782 , \REGF/pbmemout1/n6033 , 
        \REGF/pbmemout1/n6120 , \REGF/pbmemout1/n6293 , \REGF/pbmemout1/n6303 , 
        \REGF/pbmemout1/n5950 , \REGF/pbmemout1/n6324 , \REGF/pbmemout1/n5977 , 
        \REGF/pbmemout1/n6014 , \REGF/pbmemout1/n6184 , \REGF/pbmemout1/n5740 , 
        \REGF/pbmemout1/n5802 , \REGF/pbmemout1/n6128 , \REGF/pbmemout1/n6218 , 
        \REGF/pbmemout1/n5992 , \REGF/pbmemout1/n6251 , \REGF/pbmemout1/n5767 , 
        \REGF/pbmemout1/n6161 , \REGF/pbmemout1/n5825 , \REGF/pbmemout1/n6146 , 
        \REGF/pbmemout1/n6276 , \REGF/pbmemout1/n5889 , \REGF/pbmemout1/n5919 , 
        \REGF/pbmemout1/n5925 , \REGF/pbmemout1/n6376 , \REGF/pbmemout1/n6046 , 
        \REGF/pbmemout1/n6061 , \REGF/pbmemout1/n5892 , \REGF/pbmemout1/n5902 , 
        \REGF/pbmemout1/n6351 , \REGF/pbmemout1/n5682 , \REGF/pbmemout1/n5712 , 
        \REGF/pbmemout1/n5735 , \REGF/pbmemout1/n5819 , \REGF/pbmemout1/n5989 , 
        \REGF/pbmemout1/n6084 , \REGF/pbmemout1/n6114 , \REGF/pbmemout1/n5850 , 
        \REGF/pbmemout1/n6224 , \REGF/pbmemout1/n5877 , \REGF/pbmemout1/n6203 , 
        \REGF/pbmemout1/n6133 , \REGF/pbmemout1/n5799 , \REGF/pbmemout1/n6288 , 
        \REGF/pbmemout1/n6318 , \REGF/pbmemout1/n6028 , \REGF/pbmemout1/n5690 , 
        \REGF/pbmemout1/n5727 , \REGF/pbmemout1/n5959 , \REGF/pbmemout1/n6096 , 
        \REGF/pbmemout1/n6106 , \REGF/pbmemout1/n5842 , \REGF/pbmemout1/n5865 , 
        \REGF/pbmemout1/n6236 , \REGF/pbmemout1/n6211 , \REGF/pbmemout1/n6381 , 
        \REGF/pbmemout1/n6121 , \REGF/pbmemout1/n5700 , \REGF/pbmemout1/n5749 , 
        \REGF/pbmemout1/n6168 , \REGF/pbmemout1/n6258 , \REGF/pbmemout1/n5937 , 
        \REGF/pbmemout1/n6364 , \REGF/pbmemout1/n6054 , \REGF/pbmemout1/n6073 , 
        \REGF/pbmemout1/n5880 , \REGF/pbmemout1/n5910 , \REGF/pbmemout1/n5752 , 
        \REGF/pbmemout1/n5810 , \REGF/pbmemout1/n6343 , \REGF/pbmemout1/n6358 , 
        \REGF/pbmemout1/n6068 , \REGF/pbmemout1/n5980 , \REGF/pbmemout1/n6243 , 
        \REGF/pbmemout1/n5775 , \REGF/pbmemout1/n6173 , \REGF/pbmemout1/n5837 , 
        \REGF/pbmemout1/n6154 , \REGF/pbmemout1/n5859 , \REGF/pbmemout1/n6264 , 
        \REGF/pbmemout1/n5790 , \REGF/pbmemout1/n6021 , \REGF/pbmemout1/n6281 , 
        \REGF/pbmemout1/n6311 , \REGF/pbmemout1/n5942 , \REGF/pbmemout1/n6336 , 
        \REGF/pbmemout1/n5965 , \REGF/pbmemout1/n6196 , \REGF/pbmemout1/n6006 , 
        \REGF/pbmemout1/n5879 , \REGF/pbmemout1/n5755 , \REGF/pbmemout1/n5772 , 
        \REGF/pbmemout1/n5797 , \REGF/pbmemout1/n6001 , \REGF/pbmemout1/n6191 , 
        \REGF/pbmemout1/n5962 , \REGF/pbmemout1/n6331 , \REGF/pbmemout1/n5945 , 
        \REGF/pbmemout1/n6286 , \REGF/pbmemout1/n6316 , \REGF/pbmemout1/n5830 , 
        \REGF/pbmemout1/n6026 , \REGF/pbmemout1/n6378 , \REGF/pbmemout1/n6048 , 
        \REGF/pbmemout1/n6263 , \REGF/pbmemout1/n6153 , \REGF/pbmemout1/n6174 , 
        \REGF/pbmemout1/n5769 , \REGF/pbmemout1/n5817 , \REGF/pbmemout1/n6244 , 
        \REGF/pbmemout1/n5987 , \REGF/pbmemout1/n6148 , \REGF/pbmemout1/n6278 , 
        \REGF/pbmemout1/n6344 , \REGF/pbmemout1/n5887 , \REGF/pbmemout1/n5917 , 
        \REGF/pbmemout1/n6074 , \REGF/pbmemout1/n6053 , \REGF/pbmemout1/n5930 , 
        \REGF/pbmemout1/n6363 , \REGF/pbmemout1/n5979 , \REGF/pbmemout1/n5697 , 
        \REGF/pbmemout1/n5707 , \REGF/pbmemout1/n5845 , \REGF/pbmemout1/n6126 , 
        \REGF/pbmemout1/n5862 , \REGF/pbmemout1/n6216 , \REGF/pbmemout1/n5685 , 
        \REGF/pbmemout1/n5720 , \REGF/pbmemout1/n6231 , \REGF/pbmemout1/n6091 , 
        \REGF/pbmemout1/n6101 , \REGF/pbmemout1/n5715 , \REGF/pbmemout1/n5732 , 
        \REGF/pbmemout1/n5857 , \REGF/pbmemout1/n6134 , \REGF/pbmemout1/n5870 , 
        \REGF/pbmemout1/n6204 , \REGF/pbmemout1/n6223 , \REGF/pbmemout1/n6113 , 
        \REGF/pbmemout1/n6083 , \REGF/pbmemout1/n6338 , \REGF/pbmemout1/n6008 , 
        \REGF/pbmemout1/n6198 , \REGF/pbmemout1/n6356 , \REGF/pbmemout1/n5895 , 
        \REGF/pbmemout1/n5905 , \REGF/pbmemout1/n6066 , \REGF/pbmemout1/n6041 , 
        \REGF/pbmemout1/n6371 , \REGF/pbmemout1/n5922 , \REGF/pbmemout1/n5822 , 
        \REGF/pbmemout1/n5839 , \REGF/pbmemout1/n6271 , \REGF/pbmemout1/n6141 , 
        \REGF/pbmemout1/n5747 , \REGF/pbmemout1/n5760 , \REGF/pbmemout1/n6166 , 
        \REGF/pbmemout1/n5805 , \REGF/pbmemout1/n6256 , \REGF/pbmemout1/n5995 , 
        \REGF/pbmemout1/n5939 , \REGF/pbmemout1/n5729 , \REGF/pbmemout1/n5785 , 
        \REGF/pbmemout1/n6013 , \REGF/pbmemout1/n6183 , \REGF/pbmemout1/n5970 , 
        \REGF/pbmemout1/n6323 , \REGF/pbmemout1/n5957 , \REGF/pbmemout1/n6294 , 
        \REGF/pbmemout1/n6304 , \REGF/pbmemout1/n6034 , \REGF/pbmemout1/n6098 , 
        \REGF/pbmemout1/n6108 , \REGF/pbmemout1/n6238 , 
        \REGF/pbmemff11/RO_DPR28B227[6] , \REGF/pbmemff11/n5133 , 
        \REGF/pbmemff11/RO_INDY389[20] , \REGF/pbmemff11/RO_INDY389[13] , 
        \REGF/pbmemff11/n5114 , \REGF/pbmemff11/RO_INDW309[10] , 
        \REGF/pbmemff11/RO_INDY389[7] , \REGF/pbmemff11/RO_INDW309[23] , 
        \REGF/pbmemff11/RO_INDW309[19] , \REGF/pbmemff11/RO_ACC147[14] , 
        \REGF/pbmemff11/RO_ACC147[27] , \REGF/pbmemff11/n5128 , 
        \REGF/pbmemff11/RO_INDY389[29] , \REGF/pbmemff11/RO_INDY389[30] , 
        \REGF/pbmemff11/RO_ACC147[19] , \REGF/pbmemff11/RO_INDW309[14] , 
        \REGF/pbmemff11/RO_INDY389[3] , \REGF/pbmemff11/RO_INDW309[27] , 
        \REGF/pbmemff11/RO_DPR28B227[2] , \REGF/pbmemff11/RO_INDY389[24] , 
        \REGF/pbmemff11/RO_INDY389[17] , \REGF/pbmemff11/RO_ACC147[23] , 
        \REGF/pbmemff11/n5096 , \REGF/pbmemff11/RO_ACC147[10] , 
        \REGF/pbmemff11/n5106 , \REGF/pbmemff11/n5121 , 
        \REGF/pbmemff11/RO_ACC147[12] , \REGF/pbmemff11/RO_ACC147[21] , 
        \REGF/pbmemff11/n5091 , \REGF/pbmemff11/n5101 , \REGF/pbmemff11/n5126 , 
        \REGF/pbmemff11/n_1556 , \REGF/pbmemff11/RO_INDY389[8] , 
        \REGF/pbmemff11/RO_INDZ429[6] , \REGF/pbmemff11/RO_DPR28B227[9] , 
        \REGF/pbmemff11/RO_DPR28B227[0] , \REGF/pbmemff11/RO_INDY389[15] , 
        \REGF/pbmemff11/RO_INDY389[26] , \REGF/pbmemff11/RO_ACC147[28] , 
        \REGF/pbmemff11/RO_ACC147[31] , \REGF/pbmemff11/RO_INDW309[16] , 
        \REGF/pbmemff11/RO_INDY389[1] , \REGF/pbmemff11/RO_INDW309[25] , 
        \REGF/pbmemff11/RO_INDY389[18] , \REGF/pbmemff11/n5098 , 
        \REGF/pbmemff11/n5108 , \REGF/pbmemff11/RO_INDW309[28] , 
        \REGF/pbmemff11/RO_INDW309[31] , \REGF/pbmemff11/n5141 , 
        \REGF/pbmemff11/RO_ACC147[25] , \REGF/pbmemff11/RO_ACC147[16] , 
        \REGF/pbmemff11/RO_INDW309[12] , \REGF/pbmemff11/RO_INDY389[5] , 
        \REGF/pbmemff11/RO_INDW309[21] , \REGF/pbmemff11/RO_DPR28B227[4] , 
        \REGF/pbmemff11/n5113 , \REGF/pbmemff11/RO_INDY389[11] , 
        \REGF/pbmemff11/RO_INDY389[22] , \REGF/pbmemff11/n5134 , 
        \REGF/pbmemff11/n5643 , \REGF/pbmemff11/n_452 , 
        \REGF/pbmemff11/RO_SPR28B268[6] , \REGF/pbmemff11/RO_DPR28B227[15] , 
        \REGF/pbmemff11/RO_DPR28B227[26] , \REGF/pbmemff11/RO_INDW309[1] , 
        \REGF/pbmemff11/RO_ACC147[5] , \REGF/pbmemff11/RO_EACC187[11] , 
        \REGF/pbmemff11/RO_INDX349[29] , \REGF/pbmemff11/RO_INDX349[30] , 
        \REGF/pbmemff11/RO_INDZ429[29] , \REGF/pbmemff11/RO_INDZ429[30] , 
        \REGF/pbmemff11/RO_EACC187[22] , \REGF/pbmemff11/RO_EACC187[7] , 
        \REGF/pbmemff11/RO_STAT5BP[3] , \REGF/pbmemff11/RO_SPR28B268[14] , 
        \REGF/pbmemff11/RO_SPR28B268[27] , \REGF/pbmemff11/RO_INDZ429[13] , 
        \REGF/pbmemff11/RO_EACC187[18] , \REGF/pbmemff11/RO_INDZ429[20] , 
        \REGF/pbmemff11/RO_INDX349[13] , \REGF/pbmemff11/RO_INDX349[20] , 
        \REGF/pbmemff11/n5090 , \REGF/pbmemff11/n5100 , 
        \REGF/pbmemff11/RO_INDW309[8] , \REGF/pbmemff11/n5112 , 
        \REGF/pbmemff11/n5127 , \REGF/pbmemff11/RO_INDX349[3] , 
        \REGF/pbmemff11/RO_EACC187[15] , \REGF/pbmemff11/RO_EACC187[26] , 
        \REGF/pbmemff11/RO_DPR28B227[11] , \REGF/pbmemff11/RO_DPR28B227[22] , 
        \REGF/pbmemff11/RO_ACC147[8] , \REGF/pbmemff11/n5135 , 
        \REGF/pbmemff11/RO_SPR28B268[19] , \REGF/pbmemff11/RO_INDW309[5] , 
        \REGF/pbmemff11/RO_SPR28B268[2] , \REGF/pbmemff11/RO_DPR28B227[18] , 
        \REGF/pbmemff11/RO_INDX349[7] , \REGF/pbmemff11/n5140 , 
        \REGF/pbmemff11/RO_INDZ429[2] , \REGF/pbmemff11/RO_INDX349[24] , 
        \REGF/pbmemff11/RO_INDX349[17] , \REGF/pbmemff11/n5099 , 
        \REGF/pbmemff11/RO_EACC187[3] , \REGF/pbmemff11/RO_SPR28B268[23] , 
        \REGF/pbmemff11/RO_INDZ429[17] , \REGF/pbmemff11/RO_INDZ429[24] , 
        \REGF/pbmemff11/RO_SPR28B268[10] , \REGF/pbmemff11/RO_ACC147[1] , 
        \REGF/pbmemff11/n5109 , \REGF/pbmemff11/RO_INDX349[15] , 
        \REGF/pbmemff11/RO_INDX349[26] , \REGF/pbmemff11/RO_INDZ429[15] , 
        \REGF/pbmemff11/RO_ACC147[3] , \REGF/pbmemff11/RO_EACC187[1] , 
        \REGF/pbmemff11/RO_INDZ429[26] , \REGF/pbmemff11/RO_SPR28B268[12] , 
        \REGF/pbmemff11/RO_SPR28B268[21] , \REGF/pbmemff11/n5129 , 
        \REGF/pbmemff11/RO_INDX349[5] , \REGF/pbmemff11/RO_INDZ429[0] , 
        \REGF/pbmemff11/RO_SPR28B268[9] , \REGF/pbmemff11/RO_DPR28B227[13] , 
        \REGF/pbmemff11/RO_DPR28B227[20] , \REGF/pbmemff11/RO_INDW309[7] , 
        \REGF/pbmemff11/RO_SPR28B268[0] , \REGF/pbmemff11/RO_INDZ429[5] , 
        \REGF/pbmemff11/n5132 , \REGF/pbmemff11/RO_EACC187[17] , 
        \REGF/pbmemff11/RO_INDZ429[9] , \REGF/pbmemff11/RO_EACC187[24] , 
        \REGF/pbmemff11/n5115 , \REGF/pbmemff11/RO_EACC187[8] , 
        \REGF/pbmemff11/n_4044 , \REGF/pbmemff11/RO_INDZ429[4] , 
        \REGF/pbmemff11/RO_INDX349[22] , \REGF/pbmemff11/n5097 , 
        \REGF/pbmemff11/n5120 , \REGF/pbmemff11/RO_INDX349[1] , 
        \REGF/pbmemff11/RO_ACC147[7] , \REGF/pbmemff11/n5107 , 
        \REGF/pbmemff11/RO_STAT5BP[1] , \REGF/pbmemff11/RO_EACC187[5] , 
        \REGF/pbmemff11/RO_SPR28B268[25] , \REGF/pbmemff11/RO_SPR28B268[16] , 
        \REGF/pbmemff11/RO_EACC187[29] , \REGF/pbmemff11/RO_EACC187[30] , 
        \REGF/pbmemff11/RO_INDZ429[11] , \REGF/pbmemff11/RO_INDZ429[22] , 
        \REGF/pbmemff11/RO_EACC187[13] , \REGF/pbmemff11/RO_INDX349[11] , 
        \REGF/pbmemff11/RO_INDX349[18] , \REGF/pbmemff11/RO_EACC187[20] , 
        \REGF/pbmemff11/RO_INDZ429[18] , \REGF/pbmemff11/RO_SPR28B268[4] , 
        \REGF/pbmemff11/RO_DPR28B227[17] , \REGF/pbmemff11/RO_DPR28B227[24] , 
        \REGF/pbmemff11/RO_INDX349[8] , \REGF/pbmemff11/RO_INDW309[3] , 
        \REGF/pbmemff11/n5087 , \REGF/pbmemff11/n5117 , 
        \REGF/pbmemff11/RO_ACC147[6] , \REGF/pbmemff11/n5130 , 
        \REGF/pbmemff11/RO_INDX349[0] , \REGF/pbmemff11/RO_EACC187[4] , 
        \REGF/pbmemff11/RO_SPR28B268[17] , \REGF/pbmemff11/RO_SPR28B268[24] , 
        \REGF/pbmemff11/RO_INDX349[23] , \REGF/pbmemff11/RO_INDX349[10] , 
        \REGF/pbmemff11/RO_EACC187[12] , \REGF/pbmemff11/RO_EACC187[28] , 
        \REGF/pbmemff11/RO_INDZ429[10] , \REGF/pbmemff11/RO_EACC187[31] , 
        \REGF/pbmemff11/RO_INDZ429[23] , \REGF/pbmemff11/RO_EACC187[21] , 
        \REGF/pbmemff11/RO_INDX349[19] , \REGF/pbmemff11/RO_INDZ429[19] , 
        \REGF/pbmemff11/n5145 , \REGF/pbmemff11/RO_DPR28B227[16] , 
        \REGF/pbmemff11/RO_DPR28B227[25] , \REGF/pbmemff11/RO_INDW309[2] , 
        \REGF/pbmemff11/RO_SPR28B268[5] , \REGF/pbmemff11/RO_INDX349[9] , 
        \REGF/pbmemff11/RO_INDZ429[14] , \REGF/pbmemff11/RO_INDZ429[27] , 
        \REGF/pbmemff11/RO_INDX349[14] , \REGF/pbmemff11/RO_INDX349[27] , 
        \REGF/pbmemff11/RO_ACC147[2] , \REGF/pbmemff11/n5139 , 
        \REGF/pbmemff11/RO_EACC187[0] , \REGF/pbmemff11/RO_SPR28B268[20] , 
        \REGF/pbmemff11/RO_SPR28B268[13] , \REGF/pbmemff11/RO_INDX349[4] , 
        \REGF/pbmemff11/RO_SPR28B268[8] , \REGF/pbmemff11/RO_INDZ429[1] , 
        \REGF/pbmemff11/RO_DPR28B227[12] , \REGF/pbmemff11/RO_DPR28B227[21] , 
        \REGF/pbmemff11/RO_INDW309[6] , \REGF/pbmemff11/RO_SPR28B268[1] , 
        \REGF/pbmemff11/RO_INDZ429[8] , \REGF/pbmemff11/n5095 , 
        \REGF/pbmemff11/n5105 , \REGF/pbmemff11/n5122 , 
        \REGF/pbmemff11/RO_EACC187[16] , \REGF/pbmemff11/RO_EACC187[25] , 
        \REGF/pbmemff11/RO_EACC187[9] , \REGF/pbmemff11/n5092 , 
        \REGF/pbmemff11/n5102 , \REGF/pbmemff11/n5125 , 
        \REGF/pbmemff11/RO_EACC187[14] , \REGF/pbmemff11/n_3464 , 
        \REGF/pbmemff11/RO_EACC187[27] , \REGF/pbmemff11/RO_SPR28B268[18] , 
        \REGF/pbmemff11/RO_DPR28B227[10] , \REGF/pbmemff11/RO_DPR28B227[23] , 
        \REGF/pbmemff11/RO_ACC147[9] , \REGF/pbmemff11/RO_INDW309[4] , 
        \REGF/pbmemff11/RO_SPR28B268[3] , \REGF/pbmemff11/RO_DPR28B227[19] , 
        \REGF/pbmemff11/RO_INDX349[6] , \REGF/pbmemff11/RO_INDZ429[3] , 
        \REGF/pbmemff11/RO_INDX349[25] , \REGF/pbmemff11/RO_INDZ429[16] , 
        \REGF/pbmemff11/RO_INDZ429[25] , \REGF/pbmemff11/n5089 , 
        \REGF/pbmemff11/RO_ACC147[0] , \REGF/pbmemff11/RO_INDX349[16] , 
        \REGF/pbmemff11/n5119 , \REGF/pbmemff11/RO_EACC187[2] , 
        \REGF/pbmemff11/RO_SPR28B268[11] , \REGF/pbmemff11/RO_SPR28B268[22] , 
        \REGF/pbmemff11/RO_DPR28B227[14] , \REGF/pbmemff11/RO_DPR28B227[27] , 
        \REGF/pbmemff11/RO_SPR28B268[7] , \REGF/pbmemff11/RO_INDW309[0] , 
        \REGF/pbmemff11/RO_EACC187[10] , \REGF/pbmemff11/RO_EACC187[23] , 
        \REGF/pbmemff11/RO_INDZ429[31] , \REGF/pbmemff11/RO_INDZ429[28] , 
        \REGF/pbmemff11/n5142 , \REGF/pbmemff11/RO_ACC147[4] , 
        \REGF/pbmemff11/RO_EACC187[6] , \REGF/pbmemff11/RO_SPR28B268[26] , 
        \REGF/pbmemff11/RO_INDX349[28] , \REGF/pbmemff11/RO_INDX349[31] , 
        \REGF/pbmemff11/RO_SPR28B268[15] , \REGF/pbmemff11/RO_INDX349[12] , 
        \REGF/pbmemff11/RO_INDX349[21] , \REGF/pbmemff11/RO_INDZ429[12] , 
        \REGF/pbmemff11/RO_EACC187[19] , \REGF/pbmemff11/RO_INDZ429[21] , 
        \REGF/pbmemff11/RO_INDZ429[7] , \REGF/pbmemff11/n5088 , 
        \REGF/pbmemff11/n5110 , \REGF/pbmemff11/n5137 , 
        \REGF/pbmemff11/RO_INDW309[9] , \REGF/pbmemff11/RO_INDX349[2] , 
        \REGF/pbmemff11/RO_INDY389[19] , \REGF/pbmemff11/n5118 , 
        \REGF/pbmemff11/RO_ACC147[24] , \REGF/pbmemff11/RO_INDW309[29] , 
        \REGF/pbmemff11/RO_INDW309[30] , \REGF/pbmemff11/RO_ACC147[17] , 
        \REGF/pbmemff11/RO_INDY389[4] , \REGF/pbmemff11/RO_INDW309[13] , 
        \REGF/pbmemff11/RO_INDW309[20] , \REGF/pbmemff11/n5093 , 
        \REGF/pbmemff11/RO_DPR28B227[5] , \REGF/pbmemff11/n5124 , 
        \REGF/pbmemff11/RO_INDY389[23] , \REGF/pbmemff11/n5103 , 
        \REGF/pbmemff11/RO_INDY389[10] , \REGF/pbmemff11/RO_ACC147[13] , 
        \REGF/pbmemff11/RO_ACC147[20] , \REGF/pbmemff11/n5136 , 
        \REGF/pbmemff11/RO_DPR28B227[8] , \REGF/pbmemff11/n5111 , 
        \REGF/pbmemff11/RO_INDY389[9] , \REGF/pbmemff11/RO_DPR28B227[1] , 
        \REGF/pbmemff11/RO_INDY389[14] , \REGF/pbmemff11/RO_INDY389[27] , 
        \REGF/pbmemff11/n5143 , \REGF/pbmemff11/RO_ACC147[29] , 
        \REGF/pbmemff11/RO_ACC147[30] , \REGF/pbmemff11/RO_INDW309[17] , 
        \REGF/pbmemff11/n_2192 , \REGF/pbmemff11/RO_ACC147[18] , 
        \REGF/pbmemff11/RO_INDW309[24] , \REGF/pbmemff11/RO_INDY389[0] , 
        \REGF/pbmemff11/n_1032 , \REGF/pbmemff11/RO_INDY389[2] , 
        \REGF/pbmemff11/RO_INDW309[15] , \REGF/pbmemff11/RO_INDW309[26] , 
        \REGF/pbmemff11/RO_DPR28B227[3] , \REGF/pbmemff11/RO_INDY389[25] , 
        \REGF/pbmemff11/RO_INDY389[16] , \REGF/pbmemff11/n5144 , 
        \REGF/pbmemff11/RO_ACC147[22] , \REGF/pbmemff11/n5086 , 
        \REGF/pbmemff11/RO_ACC147[11] , \REGF/pbmemff11/n5094 , 
        \REGF/pbmemff11/n5104 , \REGF/pbmemff11/n5116 , \REGF/pbmemff11/n5131 , 
        \REGF/pbmemff11/RO_DPR28B227[7] , \REGF/pbmemff11/n5123 , 
        \REGF/pbmemff11/RO_INDY389[12] , \REGF/pbmemff11/RO_INDY389[21] , 
        \REGF/pbmemff11/RO_INDW309[11] , \REGF/pbmemff11/RO_ACC147[15] , 
        \REGF/pbmemff11/RO_INDW309[22] , \REGF/pbmemff11/RO_INDY389[6] , 
        \REGF/pbmemff11/RO_INDW309[18] , \REGF/pbmemff11/RO_ACC147[26] , 
        \REGF/pbmemff11/RO_INDY389[28] , \REGF/pbmemff11/RO_INDY389[31] , 
        \REGF/pbmemff11/n5138 , \MAIN/ENGIN/a_cfctl_st , \MAIN/ENGIN/n3600 , 
        \MAIN/ENGIN/b_d2_stage , \MAIN/ENGIN/b_step_end , 
        \MAIN/ENGIN/c_deocenh , \MAIN/ENGIN/status_wr4 , \MAIN/ENGIN/n3595 , 
        \MAIN/ENGIN/a_decctl_st , \MAIN/ENGIN/a_exectl_st , 
        \MAIN/ENGIN/cf_start , \MAIN/ENGIN/n3592 , \MAIN/ENGIN/status_wr3 , 
        \MAIN/ENGIN/d_d2_stage , \MAIN/ENGIN/d_step_end , \MAIN/ENGIN/n3607 , 
        \MAIN/ENGIN/D_PED4_BR , \MAIN/ENGIN/b_cf_stage , 
        \MAIN/ENGIN/c_dec_start , \MAIN/ENGIN/status_wr2 , 
        \MAIN/ENGIN/c_cfctl_st , \MAIN/ENGIN/D_INIT_STAGE , 
        \MAIN/ENGIN/d_swctl_st , \MAIN/ENGIN/n3593 , \MAIN/ENGIN/a_swctl_st , 
        \MAIN/ENGIN/a_dec_stage , \MAIN/ENGIN/b_dec_start , 
        \MAIN/ENGIN/a_deocenh , \MAIN/ENGIN/a_cf_start2 , 
        \MAIN/ENGIN/puls_exec , \MAIN/ENGIN/cf_st2_rst , 
        \MAIN/ENGIN/d_dec_start , \MAIN/ENGIN/dec_st2_rst , 
        \MAIN/ENGIN/B_PED4_BR , \MAIN/ENGIN/c_decctl_st , 
        \MAIN/ENGIN/C_INIT_STAGE , \MAIN/ENGIN/n3601 , \MAIN/ENGIN/b_swctl_st , 
        \MAIN/ENGIN/d_cf_stage , \MAIN/ENGIN/b_decctl_st , 
        \MAIN/ENGIN/d_decctl_st , \MAIN/ENGIN/n3594 , \MAIN/ENGIN/a_cf_stage , 
        \MAIN/ENGIN/A_PED4_BR , \MAIN/ENGIN/n_164 , \MAIN/ENGIN/n3603 , 
        \MAIN/ENGIN/b_deocenh , \MAIN/ENGIN/n3596 , \MAIN/ENGIN/status_wr1 , 
        \MAIN/ENGIN/n3591 , \MAIN/ENGIN/c_d2_stage , \MAIN/ENGIN/c_step_end , 
        \MAIN/ENGIN/n3604 , \MAIN/ENGIN/n3598 , \MAIN/ENGIN/b_dec_stage , 
        \MAIN/ENGIN/c_swctl_st , \MAIN/ENGIN/c_dec_stage , 
        \MAIN/ENGIN/d_cfctl_st , \MAIN/ENGIN/C_PED4_BR , 
        \MAIN/ENGIN/d_dec_stage , \MAIN/ENGIN/a_dec_start2 , 
        \MAIN/ENGIN/A_INIT_STAGE , \MAIN/ENGIN/n3599 , \MAIN/ENGIN/b_cfctl_st , 
        \MAIN/ENGIN/B_INIT_STAGE , \MAIN/ENGIN/c_cf_stage , \MAIN/ENGIN/n3602 , 
        \MAIN/ENGIN/b_exectl_st , \MAIN/ENGIN/d_exectl_st , 
        \MAIN/ENGIN/a_d2_stage , \MAIN/ENGIN/a_step_end , 
        \MAIN/ENGIN/c_exectl_st , \MAIN/ENGIN/n3597 , \MAIN/ENGIN/d_deocenh , 
        \MAIN/ENGIN/dec_start , \MAIN/ENGIN/a_dec_start , 
        \REGF/pbmemff51/n4474 , \REGF/pbmemff51/n4473 , \REGF/pbmemff51/n4469 , 
        \REGF/pbmemff51/n4472 , \REGF/pbmemff51/n4475 , \REGF/pbmemff51/n4477 , 
        \REGF/pbmemff51/n4470 , \REGF/pbmemff51/n4471 , \REGF/pbmemff51/n4476 , 
        \UPIF/CSGN/n1644 , \UPIF/CSGN/n1678 , \UPIF/CSGN/n1744 , 
        \UPIF/CSGN/n1686 , \UPIF/CSGN/n1663 , \UPIF/CSGN/n1716 , 
        \UPIF/CSGN/n1731 , \UPIF/CSGN/n1638 , \UPIF/CSGN/n1694 , 
        \UPIF/CSGN/n1704 , \UPIF/CSGN/n1723 , \UPIF/CSGN/n1656 , 
        \UPIF/CSGN/n1671 , \UPIF/CSGN/n1738 , \UPIF/CSGN/n1756 , 
        \UPIF/CSGN/n1688 , \UPIF/CSGN/n1718 , \UPIF/CSGN/n1751 , 
        \UPIF/CSGN/n1724 , \UPIF/CSGN/n1676 , \UPIF/CSGN/n1651 , 
        \UPIF/CSGN/n1681 , \UPIF/CSGN/n1693 , \UPIF/CSGN/n1736 , 
        \UPIF/CSGN/n1703 , \UPIF/CSGN/n1711 , \UPIF/CSGN/n1743 , 
        \UPIF/CSGN/n1664 , \UPIF/CSGN/n1758 , \UPIF/CSGN/n1643 , 
        \UPIF/CSGN/n1658 , \UPIF/CSGN/n1725 , \UPIF/CSGN/n1692 , 
        \UPIF/CSGN/n1702 , \UPIF/CSGN/n1650 , \UPIF/CSGN/n1677 , 
        \UPIF/CSGN/n1689 , \UPIF/CSGN/n1719 , \UPIF/CSGN/n1750 , 
        \UPIF/CSGN/n1665 , \UPIF/CSGN/n1659 , \UPIF/CSGN/n1742 , 
        \UPIF/CSGN/n1642 , \UPIF/CSGN/n1737 , \UPIF/CSGN/n1759 , 
        \UPIF/CSGN/n1710 , \UPIF/CSGN/n1680 , \UPIF/CSGN/n1687 , 
        \UPIF/CSGN/n1717 , \UPIF/CSGN/n1730 , \UPIF/CSGN/n1645 , 
        \UPIF/CSGN/n1662 , \UPIF/CSGN/n1745 , \UPIF/CSGN/n1679 , 
        \UPIF/CSGN/n1739 , \UPIF/CSGN/n1757 , \UPIF/CSGN/n1657 , 
        \UPIF/CSGN/*cell*4224/U3/CONTROL1 , \UPIF/CSGN/n1670 , 
        \UPIF/CSGN/n1639 , \UPIF/CSGN/n1705 , \UPIF/CSGN/n1695 , 
        \UPIF/CSGN/n1722 , \UPIF/CSGN/n1729 , \UPIF/CSGN/n1747 , 
        \UPIF/CSGN/n1660 , \UPIF/CSGN/n1647 , \UPIF/CSGN/n1715 , 
        \UPIF/CSGN/n1732 , \UPIF/CSGN/n1697 , \UPIF/CSGN/n1685 , 
        \UPIF/CSGN/n1720 , \UPIF/CSGN/n1707 , \UPIF/CSGN/n1672 , 
        \UPIF/CSGN/n1655 , \UPIF/CSGN/n1669 , \UPIF/CSGN/n_1054 , 
        \UPIF/CSGN/n1755 , \UPIF/CSGN/n1752 , \UPIF/CSGN/n1675 , 
        \UPIF/CSGN/n1649 , \UPIF/CSGN/n1652 , \UPIF/CSGN/n1749 , 
        \UPIF/CSGN/n1690 , \UPIF/CSGN/n1700 , \UPIF/CSGN/n1727 , 
        \UPIF/CSGN/reg_stat_h , \UPIF/CSGN/n1682 , \UPIF/CSGN/n1712 , 
        \UPIF/CSGN/n1735 , \UPIF/CSGN/n1667 , \UPIF/CSGN/n1640 , 
        \UPIF/CSGN/n1740 , \UPIF/CSGN/n1691 , \UPIF/CSGN/n1699 , 
        \UPIF/CSGN/n1709 , \UPIF/CSGN/n1701 , \UPIF/CSGN/n1726 , 
        \UPIF/CSGN/n1674 , \UPIF/CSGN/n1653 , \UPIF/CSGN/n1748 , 
        \UPIF/CSGN/n1648 , \UPIF/CSGN/n1753 , \UPIF/CSGN/n1708 , 
        \UPIF/CSGN/n1698 , \UPIF/CSGN/n_1040 , \UPIF/CSGN/n1741 , 
        \UPIF/CSGN/n1683 , \UPIF/CSGN/n1713 , \UPIF/CSGN/n1666 , 
        \UPIF/CSGN/n1641 , \UPIF/CSGN/n1714 , \UPIF/CSGN/n1734 , 
        \UPIF/CSGN/n1684 , \UPIF/CSGN/n1733 , \UPIF/CSGN/n1661 , 
        \UPIF/CSGN/n1646 , \UPIF/CSGN/n1746 , \UPIF/CSGN/n_1047 , 
        \UPIF/CSGN/n1728 , \UPIF/CSGN/n1668 , \UPIF/CSGN/n1754 , 
        \UPIF/CSGN/n1673 , \UPIF/CSGN/n1706 , \UPIF/CSGN/n1654 , 
        \UPIF/CSGN/n1721 , \UPIF/CSGN/n1696 , \CONS/phinc20_1/gg_out[2] , 
        \CONS/phinc20_1/gp_out[3] , \CONS/phinc20_1/gp_out[1] , 
        \CONS/phinc20_1/gp_out[0] , \CONS/phinc20_1/gp_out[2] , 
        \CONS/phinc20_1/gg_out[1] , \CONS/phinc20_1/gg_out[3] , 
        \CODEIF/inc19_1/gg_out[2] , \CODEIF/inc19_1/gp_out[3] , 
        \CODEIF/inc19_1/gp_out[1] , \CODEIF/inc19_1/gp_out[0] , 
        \CODEIF/inc19_1/n3764 , \CODEIF/inc19_1/n3763 , 
        \CODEIF/inc19_1/gp_out[2] , \CODEIF/inc19_1/gg_out[1] , 
        \CODEIF/inc19_1/gg_out[3] , \UPIF/RCTL/reg_file_h , \UPIF/RCTL/n1029 , 
        \UPIF/RCTL/n1032 , \UPIF/RCTL/n1035 , \UPIF/RCTL/n1040 , 
        \UPIF/RCTL/n1027 , \UPIF/RCTL/reg_eoc , \UPIF/RCTL/n1023 , 
        \UPIF/RCTL/nrt[0] , \UPIF/RCTL/n1026 , \UPIF/RCTL/irt[2] , 
        \UPIF/RCTL/n1041 , \UPIF/RCTL/n1034 , \UPIF/RCTL/irt[0] , 
        \UPIF/RCTL/n1033 , \UPIF/RCTL/nrt[2] , \UPIF/RCTL/n1028 , 
        \UPIF/RCTL/n1038 , \UPIF/RCTL/irt[1] , \UPIF/RCTL/nrt[3] , 
        \UPIF/RCTL/n_837 , \UPIF/RCTL/n1024 , \UPIF/RCTL/n1031 , 
        \UPIF/RCTL/n_839 , \UPIF/RCTL/n1036 , \UPIF/RCTL/nrt[1] , 
        \UPIF/RCTL/irt[3] , \UPIF/RCTL/n1037 , \UPIF/RCTL/n1042 , 
        \UPIF/RCTL/*cell*4328/U25/CONTROL2 , \UPIF/RCTL/n1025 , 
        \UPIF/RCTL/n_831 , \UPIF/RCTL/n1039 , \UPIF/RCTL/n1030 , 
        \CONS/lte_124/n72 , \CONS/lte_124/n287 , \CONS/lte_124/n279 , 
        \CONS/lte_124/n69 , \CONS/lte_124/n295 , \CONS/lte_124/n305 , 
        \CONS/lte_124/n67 , \CONS/lte_124/n292 , \CONS/lte_124/n302 , 
        \CONS/lte_124/n289 , \CONS/lte_124/n280 , \CONS/lte_124/n310 , 
        \CONS/lte_124/n288 , \CONS/lte_124/n63 , \CONS/lte_124/n66 , 
        \CONS/lte_124/n293 , \CONS/lte_124/n303 , \CONS/lte_124/n281 , 
        \CONS/lte_124/n68 , \CONS/lte_124/n73 , \CONS/lte_124/n278 , 
        \CONS/lte_124/n286 , \CONS/lte_124/n294 , \CONS/lte_124/n304 , 
        \CONS/lte_124/n71 , \CONS/lte_124/n284 , \CONS/lte_124/n64 , 
        \CONS/lte_124/n296 , \CONS/lte_124/n306 , \CONS/lte_124/n65 , 
        \CONS/lte_124/n291 , \CONS/lte_124/n301 , \CONS/lte_124/n298 , 
        \CONS/lte_124/n308 , \CONS/lte_124/n283 , \CONS/lte_124/n290 , 
        \CONS/lte_124/n300 , \CONS/lte_124/n282 , \CONS/lte_124/n299 , 
        \CONS/lte_124/n309 , \CONS/lte_124/n70 , \CONS/lte_124/n285 , 
        \CONS/lte_124/n297 , \CONS/lte_124/n307 , \SADR/ADRFF/n9119 , 
        \SADR/ADRFF/n9122 , \SADR/ADRFF/n9120 , \SADR/ADRFF/n9121 , 
        \SADR/ADRFF/n9123 , \SADR/ADRFF/n9124 , \REGF/pbmemff31/n5649 , 
        \REGF/pbmemff31/DO_SACONS , \REGF/pbmemff31/*cell*5410/U2/CONTROL1 , 
        \REGF/pbmemff31/RO_EST13B291[1] , \REGF/pbmemff31/n6437 , 
        \REGF/pbmemff31/n5650 , \REGF/pbmemff31/n5651 , 
        \REGF/pbmemff31/RO_PSTA3B212[1] , 
        \REGF/pbmemff31/*cell*5410/U10/CONTROL1 , 
        \REGF/pbmemff31/RO_PSTA3B212[0] , \REGF/pbmemff31/n_729 , 
        \REGF/pbmemff31/n5648 , \REGF/pbmemff31/RO_EST13B291[2] , 
        \REGF/pbmemff31/n5652 , \REGF/pbmemff31/n5647 , 
        \REGF/pbmemff31/RO_EST13B291[0] , 
        \REGF/pbmemff31/*cell*5410/U9/CONTROL1 , \SAEXE/SRCRD/nrst[0] , 
        \SAEXE/SRCRD/n93 , \SAEXE/SRCRD/erst[0] , \ALUSHT/ALU/pkdecout[31] , 
        \ALUSHT/ALU/pkdecout[28] , \ALUSHT/ALU/pkdecout[27] , 
        \ALUSHT/ALU/pkdecout[9] , \ALUSHT/ALU/pkaddsum[9] , 
        \ALUSHT/ALU/pkaddsum[0] , \ALUSHT/ALU/pkincout[26] , 
        \ALUSHT/ALU/pkincout[15] , \ALUSHT/ALU/n2180 , \ALUSHT/ALU/n2010 , 
        \ALUSHT/ALU/n1868 , \ALUSHT/ALU/n1954 , \ALUSHT/ALU/n1973 , 
        \ALUSHT/ALU/n2037 , \ALUSHT/ALU/pkaddina[26] , \ALUSHT/ALU/intb[22] , 
        \ALUSHT/ALU/intb[18] , \ALUSHT/ALU/n1806 , \ALUSHT/ALU/n1821 , 
        \ALUSHT/ALU/n1996 , \ALUSHT/ALU/n2142 , \ALUSHT/ALU/n2272 , 
        \ALUSHT/ALU/n2165 , \ALUSHT/ALU/n2255 , \ALUSHT/ALU/n2059 , 
        \ALUSHT/ALU/n2042 , \ALUSHT/ALU/n1896 , \ALUSHT/ALU/n1906 , 
        \ALUSHT/ALU/n2065 , \ALUSHT/ALU/n1921 , \ALUSHT/ALU/n2159 , 
        \ALUSHT/ALU/pkaddina[15] , \ALUSHT/ALU/pkincin[2] , \ALUSHT/ALU/n2137 , 
        \ALUSHT/ALU/n2269 , \ALUSHT/ALU/n2080 , \ALUSHT/ALU/n1854 , 
        \ALUSHT/ALU/n2207 , \ALUSHT/ALU/n1873 , \ALUSHT/ALU/n2220 , 
        \ALUSHT/ALU/n2110 , \ALUSHT/ALU/pkaddsum[4] , 
        \ALUSHT/ALU/pkaddina[18] , \ALUSHT/ALU/pkcmpinb[31] , 
        \ALUSHT/ALU/n1968 , \ALUSHT/ALU/n1846 , \ALUSHT/ALU/n2019 , 
        \ALUSHT/ALU/n2125 , \ALUSHT/ALU/n2189 , \ALUSHT/ALU/n2215 , 
        \ALUSHT/ALU/n1861 , \ALUSHT/ALU/n2232 , \ALUSHT/ALU/n2092 , 
        \ALUSHT/ALU/n2102 , \ALUSHT/ALU/pkaddina[22] , 
        \ALUSHT/ALU/pkincout[22] , \ALUSHT/ALU/pkincout[11] , 
        \ALUSHT/ALU/n2077 , \ALUSHT/ALU/n1828 , \ALUSHT/ALU/n1884 , 
        \ALUSHT/ALU/n1914 , \ALUSHT/ALU/n1933 , \ALUSHT/ALU/n2050 , 
        \ALUSHT/ALU/pkincout[18] , \ALUSHT/ALU/n1833 , \ALUSHT/ALU/n1928 , 
        \ALUSHT/ALU/n2260 , \ALUSHT/ALU/pkincin[6] , \ALUSHT/ALU/n2247 , 
        \ALUSHT/ALU/n1814 , \ALUSHT/ALU/n2150 , \ALUSHT/ALU/n2177 , 
        \ALUSHT/ALU/n1984 , \ALUSHT/ALU/pkaddina[20] , 
        \ALUSHT/ALU/pkaddina[11] , \ALUSHT/ALU/n2119 , \ALUSHT/ALU/n2089 , 
        \ALUSHT/ALU/n2229 , \ALUSHT/ALU/intb[26] , \ALUSHT/ALU/n2002 , 
        \ALUSHT/ALU/n2192 , \ALUSHT/ALU/n1946 , \ALUSHT/ALU/n1961 , 
        \ALUSHT/ALU/n2285 , \ALUSHT/ALU/n2025 , \ALUSHT/ALU/pkincin[4] , 
        \ALUSHT/ALU/n2139 , \ALUSHT/ALU/pkaddina[13] , \ALUSHT/ALU/intb[24] , 
        \ALUSHT/ALU/n2209 , \ALUSHT/ALU/intb[17] , \ALUSHT/ALU/pkincout[30] , 
        \ALUSHT/ALU/pkincout[29] , \ALUSHT/ALU/n2022 , \ALUSHT/ALU/n1908 , 
        \ALUSHT/ALU/n1941 , \ALUSHT/ALU/n1966 , \ALUSHT/ALU/n2282 , 
        \ALUSHT/ALU/n2005 , \ALUSHT/ALU/n2195 , \ALUSHT/ALU/n1898 , 
        \ALUSHT/ALU/n2240 , \ALUSHT/ALU/pkdecin[12] , \ALUSHT/ALU/pkaddsum[6] , 
        \ALUSHT/ALU/n2157 , \ALUSHT/ALU/n2170 , \ALUSHT/ALU/n1813 , 
        \ALUSHT/ALU/n1983 , \ALUSHT/ALU/n2267 , \ALUSHT/ALU/n1834 , 
        \ALUSHT/ALU/pkaddsum[2] , \ALUSHT/ALU/pkaddina[30] , 
        \ALUSHT/ALU/pkincout[20] , \ALUSHT/ALU/pkincout[13] , 
        \ALUSHT/ALU/n1808 , \ALUSHT/ALU/n1998 , \ALUSHT/ALU/n1934 , 
        \ALUSHT/ALU/n2057 , \ALUSHT/ALU/n2070 , \ALUSHT/ALU/n1883 , 
        \ALUSHT/ALU/n1913 , \ALUSHT/ALU/pkaddina[29] , 
        \ALUSHT/ALU/pkaddina[24] , \ALUSHT/ALU/intb[20] , \ALUSHT/ALU/n2045 , 
        \ALUSHT/ALU/n2095 , \ALUSHT/ALU/n2039 , \ALUSHT/ALU/n2105 , 
        \ALUSHT/ALU/n1841 , \ALUSHT/ALU/n1866 , \ALUSHT/ALU/n2235 , 
        \ALUSHT/ALU/n1853 , \ALUSHT/ALU/n1874 , \ALUSHT/ALU/n2087 , 
        \ALUSHT/ALU/n2122 , \ALUSHT/ALU/n2212 , \ALUSHT/ALU/n2117 , 
        \ALUSHT/ALU/n2227 , \ALUSHT/ALU/n1926 , \ALUSHT/ALU/n1948 , 
        \ALUSHT/ALU/n2130 , \ALUSHT/ALU/n2200 , \ALUSHT/ALU/n1891 , 
        \ALUSHT/ALU/n2062 , \ALUSHT/ALU/n1901 , \ALUSHT/ALU/pkaddina[17] , 
        \ALUSHT/ALU/pkincin[0] , \ALUSHT/ALU/n2179 , \ALUSHT/ALU/n2249 , 
        \ALUSHT/ALU/intb[30] , \ALUSHT/ALU/intb[29] , \ALUSHT/ALU/n2145 , 
        \ALUSHT/ALU/n1991 , \ALUSHT/ALU/n2252 , \ALUSHT/ALU/n2162 , 
        \ALUSHT/ALU/n1826 , \ALUSHT/ALU/n2275 , \ALUSHT/ALU/pkincin[9] , 
        \ALUSHT/ALU/n2079 , \ALUSHT/ALU/pkincout[24] , 
        \ALUSHT/ALU/pkincout[17] , \ALUSHT/ALU/n2030 , \ALUSHT/ALU/n1953 , 
        \ALUSHT/ALU/n2290 , \ALUSHT/ALU/n1974 , \ALUSHT/ALU/n1848 , 
        \ALUSHT/ALU/n2017 , \ALUSHT/ALU/n2187 , \ALUSHT/ALU/pkaddina[7] , 
        \ALUSHT/ALU/pkaddinb[21] , \ALUSHT/ALU/pkaddinb[12] , 
        \ALUSHT/ALU/inta[25] , \ALUSHT/ALU/inta[16] , \ALUSHT/ALU/n2094 , 
        \ALUSHT/ALU/n2038 , \ALUSHT/ALU/n2104 , \ALUSHT/ALU/pkaddinb[4] , 
        \ALUSHT/ALU/n2213 , \ALUSHT/ALU/n1867 , \ALUSHT/ALU/n2234 , 
        \ALUSHT/ALU/n1840 , \ALUSHT/ALU/n2123 , \ALUSHT/ALU/pkdecout[0] , 
        \ALUSHT/ALU/pkdecin[21] , \ALUSHT/ALU/pkdecin[1] , 
        \ALUSHT/ALU/pkaddsum[17] , \ALUSHT/ALU/n1809 , \ALUSHT/ALU/n1999 , 
        \ALUSHT/ALU/pkincin[23] , \ALUSHT/ALU/n1935 , 
        \ALUSHT/ALU/pkaddsum[24] , \ALUSHT/ALU/pkincin[10] , 
        \ALUSHT/ALU/n1909 , \ALUSHT/ALU/n1882 , \ALUSHT/ALU/n2056 , 
        \ALUSHT/ALU/n2071 , \ALUSHT/ALU/n1899 , \ALUSHT/ALU/n1912 , 
        \ALUSHT/ALU/pkdecin[31] , \ALUSHT/ALU/pkdecin[28] , 
        \ALUSHT/ALU/pkdecin[8] , \ALUSHT/ALU/pkincout[2] , 
        \ALUSHT/ALU/pkincin[19] , \ALUSHT/ALU/n1812 , \ALUSHT/ALU/n1982 , 
        \ALUSHT/ALU/n2171 , \ALUSHT/ALU/n2241 , \ALUSHT/ALU/n1835 , 
        \ALUSHT/ALU/n2156 , \ALUSHT/ALU/n2266 , \ALUSHT/ALU/pkdecout[23] , 
        \ALUSHT/ALU/pkdecout[19] , \ALUSHT/ALU/pkdecout[14] , 
        \ALUSHT/ALU/n2138 , \ALUSHT/ALU/pkdecin[25] , \ALUSHT/ALU/pkdecin[16] , 
        \ALUSHT/ALU/pkdecin[5] , \ALUSHT/ALU/pkaddinb[31] , \ALUSHT/ALU/n2208 , 
        \ALUSHT/ALU/pkaddinb[28] , \ALUSHT/ALU/n1940 , \ALUSHT/ALU/n2023 , 
        \ALUSHT/ALU/n2283 , \ALUSHT/ALU/n1952 , \ALUSHT/ALU/n1967 , 
        \ALUSHT/ALU/n2004 , \ALUSHT/ALU/n2031 , \ALUSHT/ALU/n2194 , 
        \ALUSHT/ALU/n2291 , \ALUSHT/ALU/pkaddsum[20] , 
        \ALUSHT/ALU/pkaddsum[13] , \ALUSHT/ALU/pkincin[27] , 
        \ALUSHT/ALU/n1975 , \ALUSHT/ALU/pkincin[14] , \ALUSHT/ALU/n2016 , 
        \ALUSHT/ALU/n2186 , \ALUSHT/ALU/n1849 , \ALUSHT/ALU/pkaddina[3] , 
        \ALUSHT/ALU/pkaddinb[0] , \ALUSHT/ALU/n1990 , \ALUSHT/ALU/n2163 , 
        \ALUSHT/ALU/n2253 , \ALUSHT/ALU/n2144 , \ALUSHT/ALU/n1827 , 
        \ALUSHT/ALU/n2274 , \ALUSHT/ALU/pkaddinb[25] , 
        \ALUSHT/ALU/pkaddinb[16] , \ALUSHT/ALU/inta[21] , \ALUSHT/ALU/n2078 , 
        \ALUSHT/ALU/pkaddinb[9] , \ALUSHT/ALU/n1927 , \ALUSHT/ALU/pkaddcin , 
        \ALUSHT/ALU/n2044 , \ALUSHT/ALU/inta[28] , \ALUSHT/ALU/n1890 , 
        \ALUSHT/ALU/n1900 , \ALUSHT/ALU/n2063 , \ALUSHT/ALU/n2178 , 
        \ALUSHT/ALU/pkdecout[21] , \ALUSHT/ALU/pkdecout[10] , 
        \ALUSHT/ALU/n2248 , \ALUSHT/ALU/pkdecout[6] , \ALUSHT/ALU/pkdecout[4] , 
        \ALUSHT/ALU/pkaddsum[30] , \ALUSHT/ALU/n2086 , \ALUSHT/ALU/n2116 , 
        \ALUSHT/ALU/pkaddsum[29] , \ALUSHT/ALU/pkincout[6] , 
        \ALUSHT/ALU/n2226 , \ALUSHT/ALU/n1852 , \ALUSHT/ALU/n1875 , 
        \ALUSHT/ALU/n2201 , \ALUSHT/ALU/n2131 , \ALUSHT/ALU/pkaddsum[18] , 
        \ALUSHT/ALU/n1949 , \ALUSHT/ALU/n2136 , \ALUSHT/ALU/pkincout[4] , 
        \ALUSHT/ALU/n1855 , \ALUSHT/ALU/n1872 , \ALUSHT/ALU/n2206 , 
        \ALUSHT/ALU/n2081 , \ALUSHT/ALU/n2221 , \ALUSHT/ALU/n2111 , 
        \ALUSHT/ALU/pkaddina[8] , \ALUSHT/ALU/n1897 , \ALUSHT/ALU/n1969 , 
        \ALUSHT/ALU/n1907 , \ALUSHT/ALU/n1920 , \ALUSHT/ALU/n2043 , 
        \ALUSHT/ALU/n2064 , \ALUSHT/ALU/pkdecout[12] , \ALUSHT/ALU/inta[19] , 
        \ALUSHT/ALU/n2158 , \ALUSHT/ALU/pkaddina[1] , \ALUSHT/ALU/n2164 , 
        \ALUSHT/ALU/n2143 , \ALUSHT/ALU/n1820 , \ALUSHT/ALU/n2268 , 
        \ALUSHT/ALU/n2273 , \ALUSHT/ALU/pkaddinb[2] , \ALUSHT/ALU/inta[23] , 
        \ALUSHT/ALU/n1807 , \ALUSHT/ALU/n2254 , \ALUSHT/ALU/n1997 , 
        \ALUSHT/ALU/pkdecout[30] , \ALUSHT/ALU/pkdecout[25] , 
        \ALUSHT/ALU/pkdecin[27] , \ALUSHT/ALU/pkdecin[14] , 
        \ALUSHT/ALU/pkdecin[7] , \ALUSHT/ALU/pkaddsum[11] , 
        \ALUSHT/ALU/pkaddinb[27] , \ALUSHT/ALU/pkaddinb[14] , 
        \ALUSHT/ALU/n2058 , \ALUSHT/ALU/pkincin[25] , \ALUSHT/ALU/n2181 , 
        \ALUSHT/ALU/n2011 , \ALUSHT/ALU/n1972 , \ALUSHT/ALU/n2296 , 
        \ALUSHT/ALU/n1955 , \ALUSHT/ALU/pkaddsum[22] , 
        \ALUSHT/ALU/pkincin[16] , \ALUSHT/ALU/n1869 , \ALUSHT/ALU/n2036 , 
        \ALUSHT/ALU/n2088 , \ALUSHT/ALU/n2118 , \ALUSHT/ALU/pkdecout[24] , 
        \ALUSHT/ALU/pkdecout[16] , \ALUSHT/ALU/n2228 , 
        \ALUSHT/ALU/pkdecout[2] , \ALUSHT/ALU/pkaddinb[19] , 
        \ALUSHT/ALU/n1929 , \ALUSHT/ALU/n1947 , \ALUSHT/ALU/n1960 , 
        \ALUSHT/ALU/n2003 , \ALUSHT/ALU/n2193 , \ALUSHT/ALU/n2024 , 
        \ALUSHT/ALU/n2284 , \ALUSHT/ALU/pkdecin[23] , \ALUSHT/ALU/pkdecin[19] , 
        \ALUSHT/ALU/pkdecin[10] , \ALUSHT/ALU/pkincout[0] , \ALUSHT/ALU/n2151 , 
        \ALUSHT/ALU/n1832 , \ALUSHT/ALU/n2261 , \ALUSHT/ALU/n2176 , 
        \ALUSHT/ALU/n2246 , \ALUSHT/ALU/pkincin[31] , \ALUSHT/ALU/n1815 , 
        \ALUSHT/ALU/n1985 , \ALUSHT/ALU/pkincin[28] , \ALUSHT/ALU/pkdecin[3] , 
        \ALUSHT/ALU/n1829 , \ALUSHT/ALU/pkaddsum[26] , 
        \ALUSHT/ALU/pkaddsum[15] , \ALUSHT/ALU/pkincout[9] , 
        \ALUSHT/ALU/n1885 , \ALUSHT/ALU/n1915 , \ALUSHT/ALU/pkincin[21] , 
        \ALUSHT/ALU/n2076 , \ALUSHT/ALU/pkaddina[5] , 
        \ALUSHT/ALU/pkaddinb[23] , \ALUSHT/ALU/pkaddinb[10] , 
        \ALUSHT/ALU/pkincin[12] , \ALUSHT/ALU/n1932 , \ALUSHT/ALU/n2051 , 
        \ALUSHT/ALU/pkaddinb[6] , \ALUSHT/ALU/inta[27] , \ALUSHT/ALU/n2018 , 
        \ALUSHT/ALU/n2188 , \ALUSHT/ALU/pkaddinb[18] , \ALUSHT/ALU/n2214 , 
        \ALUSHT/ALU/n1847 , \ALUSHT/ALU/n2124 , \ALUSHT/ALU/n2103 , 
        \ALUSHT/ALU/n1860 , \ALUSHT/ALU/n2233 , \ALUSHT/ALU/n2093 , 
        \ALUSHT/ALU/pkdecout[20] , \ALUSHT/ALU/pkdecout[17] , 
        \ALUSHT/ALU/n2098 , \ALUSHT/ALU/n2108 , \ALUSHT/ALU/pkdecout[7] , 
        \ALUSHT/ALU/pkdecout[3] , \ALUSHT/ALU/n2034 , \ALUSHT/ALU/n1957 , 
        \ALUSHT/ALU/n2238 , \ALUSHT/ALU/n2294 , \ALUSHT/ALU/n1970 , 
        \ALUSHT/ALU/n2013 , \ALUSHT/ALU/n2183 , \ALUSHT/ALU/pkdecin[22] , 
        \ALUSHT/ALU/pkdecin[18] , \ALUSHT/ALU/pkdecin[11] , 
        \ALUSHT/ALU/pkincout[1] , \ALUSHT/ALU/pkincin[30] , 
        \ALUSHT/ALU/pkincin[29] , \ALUSHT/ALU/n1805 , \ALUSHT/ALU/n1939 , 
        \ALUSHT/ALU/n2166 , \ALUSHT/ALU/n1995 , \ALUSHT/ALU/n2256 , 
        \ALUSHT/ALU/n1822 , \ALUSHT/ALU/n1839 , \ALUSHT/ALU/n2141 , 
        \ALUSHT/ALU/n2271 , \ALUSHT/ALU/pkdecin[2] , \ALUSHT/ALU/pkaddsum[14] , 
        \ALUSHT/ALU/pkincin[20] , \ALUSHT/ALU/n1895 , \ALUSHT/ALU/n1922 , 
        \ALUSHT/ALU/n2041 , \ALUSHT/ALU/n1905 , \ALUSHT/ALU/pkaddsum[27] , 
        \ALUSHT/ALU/pkincout[8] , \ALUSHT/ALU/pkincin[13] , 
        \ALUSHT/ALU/pkaddsum[19] , \ALUSHT/ALU/pkaddina[4] , 
        \ALUSHT/ALU/pkaddinb[22] , \ALUSHT/ALU/pkaddinb[11] , 
        \ALUSHT/ALU/inta[26] , \ALUSHT/ALU/n2066 , \ALUSHT/ALU/n2008 , 
        \ALUSHT/ALU/n2198 , \ALUSHT/ALU/n2083 , \ALUSHT/ALU/n1870 , 
        \ALUSHT/ALU/n2223 , \ALUSHT/ALU/n2113 , \ALUSHT/ALU/n2134 , 
        \ALUSHT/ALU/pkaddinb[7] , \ALUSHT/ALU/pkincout[5] , \ALUSHT/ALU/n2101 , 
        \ALUSHT/ALU/n1857 , \ALUSHT/ALU/n2204 , \ALUSHT/ALU/n1862 , 
        \ALUSHT/ALU/n2231 , \ALUSHT/ALU/n2091 , \ALUSHT/ALU/n2126 , 
        \ALUSHT/ALU/n2216 , \ALUSHT/ALU/n1845 , \ALUSHT/ALU/n1979 , 
        \ALUSHT/ALU/pkaddina[9] , \ALUSHT/ALU/n1887 , \ALUSHT/ALU/n1917 , 
        \ALUSHT/ALU/n1930 , \ALUSHT/ALU/n2053 , \ALUSHT/ALU/n2074 , 
        \ALUSHT/ALU/n2148 , \ALUSHT/ALU/pkdecout[13] , \ALUSHT/ALU/n2278 , 
        \ALUSHT/ALU/pkaddina[0] , \ALUSHT/ALU/pkaddinb[3] , 
        \ALUSHT/ALU/inta[18] , \ALUSHT/ALU/pkaddinb[26] , 
        \ALUSHT/ALU/pkaddinb[15] , \ALUSHT/ALU/n2244 , \ALUSHT/ALU/n1817 , 
        \ALUSHT/ALU/n1987 , \ALUSHT/ALU/n2174 , \ALUSHT/ALU/n2153 , 
        \ALUSHT/ALU/n1830 , \ALUSHT/ALU/n2263 , \ALUSHT/ALU/n2048 , 
        \ALUSHT/ALU/pkdecout[29] , \ALUSHT/ALU/pkdecout[26] , 
        \ALUSHT/ALU/pkdecout[22] , \ALUSHT/ALU/pkdecout[18] , 
        \ALUSHT/ALU/pkdecin[26] , \ALUSHT/ALU/pkdecin[15] , 
        \ALUSHT/ALU/pkdecin[6] , \ALUSHT/ALU/inta[22] , 
        \ALUSHT/ALU/pkaddsum[23] , \ALUSHT/ALU/pkaddsum[10] , 
        \ALUSHT/ALU/n2286 , \ALUSHT/ALU/pkincin[24] , \ALUSHT/ALU/n2026 , 
        \ALUSHT/ALU/n1945 , \ALUSHT/ALU/pkincin[17] , \ALUSHT/ALU/n1962 , 
        \ALUSHT/ALU/n2001 , \ALUSHT/ALU/n2191 , \ALUSHT/ALU/pkdecin[24] , 
        \ALUSHT/ALU/pkdecin[17] , \ALUSHT/ALU/pkdecin[4] , 
        \ALUSHT/ALU/pkaddsum[12] , \ALUSHT/ALU/pkcmpina[31] , 
        \ALUSHT/ALU/n1879 , \ALUSHT/ALU/n1965 , \ALUSHT/ALU/pkincin[26] , 
        \ALUSHT/ALU/pkaddsum[21] , \ALUSHT/ALU/pkincin[15] , 
        \ALUSHT/ALU/n2006 , \ALUSHT/ALU/n1942 , \ALUSHT/ALU/n2021 , 
        \ALUSHT/ALU/n2196 , \ALUSHT/ALU/n2281 , \ALUSHT/ALU/pkaddina[2] , 
        \ALUSHT/ALU/n1859 , \ALUSHT/ALU/n2154 , \ALUSHT/ALU/pkaddinb[24] , 
        \ALUSHT/ALU/pkaddinb[17] , \ALUSHT/ALU/pkaddinb[1] , 
        \ALUSHT/ALU/pkeqflg , \ALUSHT/ALU/n1810 , \ALUSHT/ALU/n1837 , 
        \ALUSHT/ALU/n2264 , \ALUSHT/ALU/n2243 , \ALUSHT/ALU/n1980 , 
        \ALUSHT/ALU/n2173 , \ALUSHT/ALU/pkaddinb[8] , \ALUSHT/ALU/inta[20] , 
        \ALUSHT/ALU/n2073 , \ALUSHT/ALU/n2068 , \ALUSHT/ALU/n1880 , 
        \ALUSHT/ALU/n1910 , \ALUSHT/ALU/n1937 , \ALUSHT/ALU/n2054 , 
        \ALUSHT/ALU/pkdecout[11] , \ALUSHT/ALU/inta[30] , 
        \ALUSHT/ALU/inta[29] , \ALUSHT/ALU/n2168 , \ALUSHT/ALU/pkdecout[8] , 
        \ALUSHT/ALU/pkdecout[5] , \ALUSHT/ALU/pkaddsum[31] , 
        \ALUSHT/ALU/pkaddsum[28] , \ALUSHT/ALU/n2258 , \ALUSHT/ALU/n1842 , 
        \ALUSHT/ALU/n2121 , \ALUSHT/ALU/n2211 , \ALUSHT/ALU/pkincout[7] , 
        \ALUSHT/ALU/n2096 , \ALUSHT/ALU/n1865 , \ALUSHT/ALU/n2106 , 
        \ALUSHT/ALU/n2236 , \ALUSHT/ALU/n1959 , \ALUSHT/ALU/pkdecin[20] , 
        \ALUSHT/ALU/pkdecin[13] , \ALUSHT/ALU/pkaddina[6] , 
        \ALUSHT/ALU/pkaddinb[20] , \ALUSHT/ALU/pkaddinb[13] , 
        \ALUSHT/ALU/inta[24] , \ALUSHT/ALU/inta[17] , \ALUSHT/ALU/n2288 , 
        \ALUSHT/ALU/n2028 , \ALUSHT/ALU/pkaddinb[5] , \ALUSHT/ALU/n1850 , 
        \ALUSHT/ALU/n2133 , \ALUSHT/ALU/n2203 , \ALUSHT/ALU/n2084 , 
        \ALUSHT/ALU/n2114 , \ALUSHT/ALU/n1819 , \ALUSHT/ALU/n1877 , 
        \ALUSHT/ALU/n1989 , \ALUSHT/ALU/n2224 , \ALUSHT/ALU/pkdecout[1] , 
        \ALUSHT/ALU/pkdecin[30] , \ALUSHT/ALU/pkdecin[29] , 
        \ALUSHT/ALU/pkdecin[0] , \ALUSHT/ALU/n1892 , \ALUSHT/ALU/n1902 , 
        \ALUSHT/ALU/n2061 , \ALUSHT/ALU/pkaddsum[25] , 
        \ALUSHT/ALU/pkaddsum[16] , \ALUSHT/ALU/pkincin[22] , 
        \ALUSHT/ALU/pkincin[11] , \ALUSHT/ALU/n2046 , \ALUSHT/ALU/n1925 , 
        \ALUSHT/ALU/pkdecin[9] , \ALUSHT/ALU/pkincout[3] , 
        \ALUSHT/ALU/pkincin[18] , \ALUSHT/ALU/n2146 , \ALUSHT/ALU/n1889 , 
        \ALUSHT/ALU/n1919 , \ALUSHT/ALU/n2276 , \ALUSHT/ALU/pkaddinb[30] , 
        \ALUSHT/ALU/pkaddinb[29] , \ALUSHT/ALU/n2251 , \ALUSHT/ALU/n1825 , 
        \ALUSHT/ALU/n1802 , \ALUSHT/ALU/n1992 , \ALUSHT/ALU/n2161 , 
        \ALUSHT/ALU/n2128 , \ALUSHT/ALU/pkdecout[15] , \ALUSHT/ALU/n2218 , 
        \ALUSHT/ALU/pkaddsum[8] , \ALUSHT/ALU/pkaddsum[7] , 
        \ALUSHT/ALU/pkaddsum[3] , \ALUSHT/ALU/pkaddina[25] , 
        \ALUSHT/ALU/n2014 , \ALUSHT/ALU/n1977 , \ALUSHT/ALU/n2184 , 
        \ALUSHT/ALU/n1843 , \ALUSHT/ALU/n1950 , \ALUSHT/ALU/n2033 , 
        \ALUSHT/ALU/n2210 , \ALUSHT/ALU/n2293 , \ALUSHT/ALU/n1864 , 
        \ALUSHT/ALU/n2097 , \ALUSHT/ALU/n2107 , \ALUSHT/ALU/n2120 , 
        \ALUSHT/ALU/n2237 , \ALUSHT/ALU/n1881 , \ALUSHT/ALU/n1958 , 
        \ALUSHT/ALU/n1911 , \ALUSHT/ALU/n2072 , \ALUSHT/ALU/n1936 , 
        \ALUSHT/ALU/n2055 , \ALUSHT/ALU/pkincin[1] , \ALUSHT/ALU/n2169 , 
        \ALUSHT/ALU/pkaddina[16] , \ALUSHT/ALU/intb[28] , 
        \ALUSHT/ALU/intb[21] , \ALUSHT/ALU/n2259 , \ALUSHT/ALU/n1836 , 
        \ALUSHT/ALU/n2155 , \ALUSHT/ALU/n1811 , \ALUSHT/ALU/n1981 , 
        \ALUSHT/ALU/n2265 , \ALUSHT/ALU/n2242 , \ALUSHT/ALU/n2172 , 
        \ALUSHT/ALU/pkincin[8] , \ALUSHT/ALU/n2069 , \ALUSHT/ALU/pkincout[25] , 
        \ALUSHT/ALU/pkincout[16] , \ALUSHT/ALU/n1964 , \ALUSHT/ALU/n2007 , 
        \ALUSHT/ALU/n2197 , \ALUSHT/ALU/n2020 , \ALUSHT/ALU/n2280 , 
        \ALUSHT/ALU/n1943 , \ALUSHT/ALU/pkaddina[21] , \ALUSHT/ALU/intb[25] , 
        \ALUSHT/ALU/n1858 , \ALUSHT/ALU/intb[16] , \ALUSHT/ALU/pkaddina[12] , 
        \ALUSHT/ALU/pkincin[5] , \ALUSHT/ALU/n2129 , \ALUSHT/ALU/n2219 , 
        \ALUSHT/ALU/pkincout[31] , \ALUSHT/ALU/n1824 , \ALUSHT/ALU/n1888 , 
        \ALUSHT/ALU/n1976 , \ALUSHT/ALU/n2015 , \ALUSHT/ALU/n2032 , 
        \ALUSHT/ALU/n2185 , \ALUSHT/ALU/n1951 , \ALUSHT/ALU/n2292 , 
        \ALUSHT/ALU/n1918 , \ALUSHT/ALU/n2147 , \ALUSHT/ALU/n1803 , 
        \ALUSHT/ALU/n2277 , \ALUSHT/ALU/n1993 , \ALUSHT/ALU/pkincout[28] , 
        \ALUSHT/ALU/n2250 , \ALUSHT/ALU/n1818 , \ALUSHT/ALU/n2160 , 
        \ALUSHT/ALU/n1988 , \ALUSHT/ALU/pkaddsum[5] , 
        \ALUSHT/ALU/pkaddina[31] , \ALUSHT/ALU/pkaddina[28] , 
        \ALUSHT/ALU/pkincout[21] , \ALUSHT/ALU/pkincout[12] , 
        \ALUSHT/ALU/n2060 , \ALUSHT/ALU/n1893 , \ALUSHT/ALU/n1903 , 
        \ALUSHT/ALU/n1924 , \ALUSHT/ALU/n2029 , \ALUSHT/ALU/n2047 , 
        \ALUSHT/ALU/n2289 , \ALUSHT/ALU/pkaddina[19] , \ALUSHT/ALU/n1851 , 
        \ALUSHT/ALU/n2202 , \ALUSHT/ALU/n1876 , \ALUSHT/ALU/n2085 , 
        \ALUSHT/ALU/n2132 , \ALUSHT/ALU/n2115 , \ALUSHT/ALU/n2225 , 
        \ALUSHT/ALU/n2135 , \ALUSHT/ALU/n2082 , \ALUSHT/ALU/n1871 , 
        \ALUSHT/ALU/n2009 , \ALUSHT/ALU/n2199 , \ALUSHT/ALU/n2112 , 
        \ALUSHT/ALU/n2222 , \ALUSHT/ALU/n1838 , \ALUSHT/ALU/n1856 , 
        \ALUSHT/ALU/n2205 , \ALUSHT/ALU/pkaddsum[1] , \ALUSHT/ALU/pkovf32 , 
        \ALUSHT/ALU/pkgtflg , \ALUSHT/ALU/pkincout[23] , 
        \ALUSHT/ALU/pkincout[10] , \ALUSHT/ALU/n2040 , \ALUSHT/ALU/n1894 , 
        \ALUSHT/ALU/n1904 , \ALUSHT/ALU/n1923 , \ALUSHT/ALU/n1938 , 
        \ALUSHT/ALU/n2067 , \ALUSHT/ALU/n1994 , \ALUSHT/ALU/n2167 , 
        \ALUSHT/ALU/n2257 , \ALUSHT/ALU/n1804 , \ALUSHT/ALU/n1823 , 
        \ALUSHT/ALU/n2270 , \ALUSHT/ALU/pkaddina[23] , \ALUSHT/ALU/intb[27] , 
        \ALUSHT/ALU/pkincout[19] , \ALUSHT/ALU/n2140 , \ALUSHT/ALU/n2109 , 
        \ALUSHT/ALU/n2099 , \ALUSHT/ALU/pkaddina[10] , \ALUSHT/ALU/pkincin[7] , 
        \ALUSHT/ALU/pkincout[27] , \ALUSHT/ALU/pkincout[14] , 
        \ALUSHT/ALU/n1956 , \ALUSHT/ALU/n2239 , \ALUSHT/ALU/n2035 , 
        \ALUSHT/ALU/n2295 , \ALUSHT/ALU/n1971 , \ALUSHT/ALU/n2012 , 
        \ALUSHT/ALU/n2182 , \ALUSHT/ALU/n1944 , \ALUSHT/ALU/n2000 , 
        \ALUSHT/ALU/n2027 , \ALUSHT/ALU/n2287 , \ALUSHT/ALU/n2190 , 
        \ALUSHT/ALU/n1963 , \ALUSHT/ALU/pkaddina[27] , \ALUSHT/ALU/intb[19] , 
        \ALUSHT/ALU/n2245 , \ALUSHT/ALU/n1878 , \ALUSHT/ALU/n2175 , 
        \ALUSHT/ALU/n2152 , \ALUSHT/ALU/n1816 , \ALUSHT/ALU/n1831 , 
        \ALUSHT/ALU/n1986 , \ALUSHT/ALU/n2262 , \ALUSHT/ALU/pkincin[3] , 
        \ALUSHT/ALU/n2075 , \ALUSHT/ALU/n1886 , \ALUSHT/ALU/n2049 , 
        \ALUSHT/ALU/n2052 , \ALUSHT/ALU/n1931 , \ALUSHT/ALU/n1916 , 
        \ALUSHT/ALU/pkaddina[14] , \ALUSHT/ALU/n2149 , \ALUSHT/ALU/n2279 , 
        \ALUSHT/ALU/intb[23] , \ALUSHT/ALU/n1844 , \ALUSHT/ALU/n1863 , 
        \ALUSHT/ALU/n2090 , \ALUSHT/ALU/n2230 , \ALUSHT/ALU/n2100 , 
        \ALUSHT/ALU/n2127 , \ALUSHT/ALU/n1978 , \ALUSHT/ALU/n2217 , 
        \ALUSHT/SHT/n2387 , \ALUSHT/SHT/n2531 , \ALUSHT/SHT/n2601 , 
        \ALUSHT/SHT/n2791 , \ALUSHT/SHT/n2943 , \ALUSHT/SHT/n3064 , 
        \ALUSHT/SHT/n2297 , \ALUSHT/SHT/n2320 , \ALUSHT/SHT/n2307 , 
        \ALUSHT/SHT/n2486 , \ALUSHT/SHT/n2964 , \ALUSHT/SHT/n2516 , 
        \ALUSHT/SHT/n2626 , \ALUSHT/SHT/n3043 , \ALUSHT/SHT/n2858 , 
        \ALUSHT/SHT/n2397 , \ALUSHT/SHT/n2774 , \ALUSHT/SHT/n2811 , 
        \ALUSHT/SHT/n2981 , \ALUSHT/SHT/n2753 , \ALUSHT/SHT/n2463 , 
        \ALUSHT/SHT/n3081 , \ALUSHT/SHT/n3111 , \ALUSHT/SHT/n3036 , 
        \ALUSHT/SHT/n2674 , \ALUSHT/SHT/n2444 , \ALUSHT/SHT/n2836 , 
        \ALUSHT/SHT/n2544 , \ALUSHT/SHT/n2648 , \ALUSHT/SHT/n2369 , 
        \ALUSHT/SHT/n2578 , \ALUSHT/SHT/n2355 , \ALUSHT/SHT/n2936 , 
        \ALUSHT/SHT/n3011 , \ALUSHT/SHT/n2478 , \ALUSHT/SHT/n2911 , 
        \ALUSHT/SHT/n2653 , \ALUSHT/SHT/n2372 , \ALUSHT/SHT/n2563 , 
        \ALUSHT/SHT/n2881 , \ALUSHT/SHT/n2748 , \ALUSHT/SHT/n2726 , 
        \ALUSHT/SHT/n2416 , \ALUSHT/SHT/n2864 , \ALUSHT/SHT/n2404 , 
        \ALUSHT/SHT/n2329 , \ALUSHT/SHT/n2701 , \ALUSHT/SHT/n2431 , 
        \ALUSHT/SHT/n2843 , \ALUSHT/SHT/n2586 , \ALUSHT/SHT/n2691 , 
        \ALUSHT/SHT/n2958 , \ALUSHT/SHT/n3058 , \ALUSHT/SHT/n2734 , 
        \ALUSHT/SHT/n2538 , \ALUSHT/SHT/n2608 , \ALUSHT/SHT/n2798 , 
        \ALUSHT/SHT/n2594 , \ALUSHT/SHT/n2385 , \ALUSHT/SHT/n2683 , 
        \ALUSHT/SHT/n2876 , \ALUSHT/SHT/n2423 , \ALUSHT/SHT/n2713 , 
        \ALUSHT/SHT/n2851 , \ALUSHT/SHT/n2918 , \ALUSHT/SHT/n2924 , 
        \ALUSHT/SHT/n2818 , \ALUSHT/SHT/n3088 , \ALUSHT/SHT/n2347 , 
        \ALUSHT/SHT/n2988 , \ALUSHT/SHT/n2556 , \ALUSHT/SHT/n3024 , 
        \ALUSHT/SHT/n2666 , \ALUSHT/SHT/n3003 , \ALUSHT/SHT/n2641 , 
        \ALUSHT/SHT/n2893 , \ALUSHT/SHT/n2360 , \ALUSHT/SHT/n2571 , 
        \ALUSHT/SHT/n2903 , \ALUSHT/SHT/n2888 , \ALUSHT/SHT/n2399 , 
        \ALUSHT/SHT/n2523 , \ALUSHT/SHT/n2438 , \ALUSHT/SHT/n2741 , 
        \ALUSHT/SHT/n3018 , \ALUSHT/SHT/n2471 , \ALUSHT/SHT/n2803 , 
        \ALUSHT/SHT/n2993 , \ALUSHT/SHT/n2698 , \ALUSHT/SHT/n2824 , 
        \ALUSHT/SHT/n2456 , \ALUSHT/SHT/n2766 , \ALUSHT/SHT/n3093 , 
        \ALUSHT/SHT/n3103 , \ALUSHT/SHT/n2708 , \ALUSHT/SHT/n2332 , 
        \ALUSHT/SHT/n2783 , \ALUSHT/SHT/n2613 , \ALUSHT/SHT/n3076 , 
        \ALUSHT/SHT/n2951 , \ALUSHT/SHT/n2634 , \ALUSHT/SHT/n2315 , 
        \ALUSHT/SHT/n2504 , \ALUSHT/SHT/n2494 , \ALUSHT/SHT/n2976 , 
        \ALUSHT/SHT/n2728 , \ALUSHT/SHT/n3051 , \ALUSHT/SHT/n2588 , 
        \ALUSHT/SHT/n2418 , \ALUSHT/SHT/n2524 , \ALUSHT/SHT/n2971 , 
        \ALUSHT/SHT/n2633 , \ALUSHT/SHT/n3056 , \ALUSHT/SHT/n2312 , 
        \ALUSHT/SHT/n2503 , \ALUSHT/SHT/n2493 , \ALUSHT/SHT/n2956 , 
        \ALUSHT/SHT/n2823 , \ALUSHT/SHT/n2335 , \ALUSHT/SHT/n2614 , 
        \ALUSHT/SHT/n3071 , \ALUSHT/SHT/n2784 , \ALUSHT/SHT/n2938 , 
        \ALUSHT/SHT/n3038 , \ALUSHT/SHT/n2451 , \ALUSHT/SHT/n2476 , 
        \ALUSHT/SHT/n2994 , \ALUSHT/SHT/n2746 , \ALUSHT/SHT/n2761 , 
        \ALUSHT/SHT/n3094 , \ALUSHT/SHT/n3104 , \ALUSHT/SHT/n2804 , 
        \ALUSHT/SHT/n2390 , \ALUSHT/SHT/n2593 , \ALUSHT/SHT/n2923 , 
        \ALUSHT/SHT/n2367 , \ALUSHT/SHT/n2904 , \ALUSHT/SHT/n2838 , 
        \ALUSHT/SHT/n2894 , \ALUSHT/SHT/n2576 , \ALUSHT/SHT/n2661 , 
        \ALUSHT/SHT/n2646 , \ALUSHT/SHT/n3023 , \ALUSHT/SHT/n3004 , 
        \ALUSHT/SHT/n2551 , \ALUSHT/SHT/n2340 , \ALUSHT/SHT/n2309 , 
        \ALUSHT/SHT/n2488 , \ALUSHT/SHT/n2299 , \ALUSHT/SHT/n2382 , 
        \ALUSHT/SHT/n2856 , \ALUSHT/SHT/n2518 , \ALUSHT/SHT/n2628 , 
        \ALUSHT/SHT/n2684 , \ALUSHT/SHT/n2714 , \ALUSHT/SHT/n2871 , 
        \ALUSHT/SHT/n2424 , \ALUSHT/SHT/n2403 , \ALUSHT/SHT/n2436 , 
        \ALUSHT/SHT/n2733 , \ALUSHT/SHT/n2696 , \ALUSHT/SHT/n2706 , 
        \ALUSHT/SHT/n2581 , \ALUSHT/SHT/n2844 , \ALUSHT/SHT/n2558 , 
        \ALUSHT/SHT/n2458 , \ALUSHT/SHT/n2654 , \ALUSHT/SHT/n2411 , 
        \ALUSHT/SHT/n2978 , \ALUSHT/SHT/n2721 , \ALUSHT/SHT/n2863 , 
        \ALUSHT/SHT/n3078 , \ALUSHT/SHT/n2375 , \ALUSHT/SHT/n2564 , 
        \ALUSHT/SHT/n2886 , \ALUSHT/SHT/n2916 , \ALUSHT/SHT/n2673 , 
        \ALUSHT/SHT/n3031 , \ALUSHT/SHT/n2931 , \ALUSHT/SHT/n2352 , 
        \ALUSHT/SHT/n2543 , \ALUSHT/SHT/n3016 , \ALUSHT/SHT/n2768 , 
        \ALUSHT/SHT/n2443 , \ALUSHT/SHT/n2831 , \ALUSHT/SHT/n2754 , 
        \ALUSHT/SHT/n2773 , \ALUSHT/SHT/n3086 , \ALUSHT/SHT/n2464 , 
        \ALUSHT/SHT/n2816 , \ALUSHT/SHT/n2986 , \ALUSHT/SHT/n2668 , 
        \ALUSHT/SHT/n2349 , \ALUSHT/SHT/n2481 , \ALUSHT/SHT/n2300 , 
        \ALUSHT/SHT/n2511 , \ALUSHT/SHT/n2621 , \ALUSHT/SHT/n3044 , 
        \ALUSHT/SHT/n2878 , \ALUSHT/SHT/n2796 , \ALUSHT/SHT/n2327 , 
        \ALUSHT/SHT/n2963 , \ALUSHT/SHT/n2536 , \ALUSHT/SHT/n2944 , 
        \ALUSHT/SHT/n3063 , \ALUSHT/SHT/n2606 , \ALUSHT/SHT/n2402 , 
        \ALUSHT/SHT/n2298 , \ALUSHT/SHT/n2519 , \ALUSHT/SHT/n2685 , 
        \ALUSHT/SHT/n2308 , \ALUSHT/SHT/n2489 , \ALUSHT/SHT/n2629 , 
        \ALUSHT/SHT/n2715 , \ALUSHT/SHT/n2857 , \ALUSHT/SHT/n2425 , 
        \ALUSHT/SHT/n2592 , \ALUSHT/SHT/n2870 , \ALUSHT/SHT/n2383 , 
        \ALUSHT/SHT/n2732 , \ALUSHT/SHT/n2922 , \ALUSHT/SHT/n2577 , 
        \ALUSHT/SHT/n2895 , \ALUSHT/SHT/n2839 , \ALUSHT/SHT/n2905 , 
        \ALUSHT/SHT/n2366 , \ALUSHT/SHT/n2647 , \ALUSHT/SHT/n3022 , 
        \ALUSHT/SHT/n2660 , \ALUSHT/SHT/n3005 , \ALUSHT/SHT/n2341 , 
        \ALUSHT/SHT/n2550 , \ALUSHT/SHT/n2939 , \ALUSHT/SHT/n2398 , 
        \ALUSHT/SHT/n2477 , \ALUSHT/SHT/n3039 , \ALUSHT/SHT/n2760 , 
        \ALUSHT/SHT/n2450 , \ALUSHT/SHT/n2822 , \ALUSHT/SHT/n3095 , 
        \ALUSHT/SHT/n3105 , \ALUSHT/SHT/n2805 , \ALUSHT/SHT/n2747 , 
        \ALUSHT/SHT/n2995 , \ALUSHT/SHT/n2729 , \ALUSHT/SHT/n2419 , 
        \ALUSHT/SHT/n2589 , \ALUSHT/SHT/n2525 , \ALUSHT/SHT/n2492 , 
        \ALUSHT/SHT/n2970 , \ALUSHT/SHT/n2632 , \ALUSHT/SHT/n3057 , 
        \ALUSHT/SHT/n2502 , \ALUSHT/SHT/n2957 , \ALUSHT/SHT/n2313 , 
        \ALUSHT/SHT/n2334 , \ALUSHT/SHT/n2480 , \ALUSHT/SHT/n2615 , 
        \ALUSHT/SHT/n2785 , \ALUSHT/SHT/n2620 , \ALUSHT/SHT/n3070 , 
        \ALUSHT/SHT/n3045 , \ALUSHT/SHT/n2945 , \ALUSHT/SHT/n2301 , 
        \ALUSHT/SHT/n2510 , \ALUSHT/SHT/n2326 , \ALUSHT/SHT/n2537 , 
        \ALUSHT/SHT/n2962 , \ALUSHT/SHT/n2879 , \ALUSHT/SHT/n2797 , 
        \ALUSHT/SHT/n2607 , \ALUSHT/SHT/n3062 , \ALUSHT/SHT/n2396 , 
        \ALUSHT/SHT/n2930 , \ALUSHT/SHT/n2669 , \ALUSHT/SHT/n2442 , 
        \ALUSHT/SHT/n2755 , \ALUSHT/SHT/n2830 , \ALUSHT/SHT/n2772 , 
        \ALUSHT/SHT/n3087 , \ALUSHT/SHT/n2817 , \ALUSHT/SHT/n2465 , 
        \ALUSHT/SHT/n2987 , \ALUSHT/SHT/n2348 , \ALUSHT/SHT/n2559 , 
        \ALUSHT/SHT/n2672 , \ALUSHT/SHT/n3030 , \ALUSHT/SHT/n2374 , 
        \ALUSHT/SHT/n2565 , \ALUSHT/SHT/n2887 , \ALUSHT/SHT/n2917 , 
        \ALUSHT/SHT/n3017 , \ALUSHT/SHT/n2655 , \ALUSHT/SHT/n2542 , 
        \ALUSHT/SHT/n2353 , \ALUSHT/SHT/n2459 , \ALUSHT/SHT/n2769 , 
        \ALUSHT/SHT/n2410 , \ALUSHT/SHT/n2437 , \ALUSHT/SHT/n2697 , 
        \ALUSHT/SHT/n2707 , \ALUSHT/SHT/n2845 , \ALUSHT/SHT/n3079 , 
        \ALUSHT/SHT/n2862 , \ALUSHT/SHT/n2391 , \ALUSHT/SHT/n2580 , 
        \ALUSHT/SHT/n2720 , \ALUSHT/SHT/n2727 , \ALUSHT/SHT/n2979 , 
        \ALUSHT/SHT/n2587 , \ALUSHT/SHT/n2865 , \ALUSHT/SHT/n2545 , 
        \ALUSHT/SHT/n2690 , \ALUSHT/SHT/n2700 , \ALUSHT/SHT/n2842 , 
        \ALUSHT/SHT/n2417 , \ALUSHT/SHT/n2430 , \ALUSHT/SHT/n2937 , 
        \ALUSHT/SHT/n2959 , \ALUSHT/SHT/n3059 , \ALUSHT/SHT/n2775 , 
        \ALUSHT/SHT/n3037 , \ALUSHT/SHT/n2354 , \ALUSHT/SHT/n2652 , 
        \ALUSHT/SHT/n2675 , \ALUSHT/SHT/n3010 , \ALUSHT/SHT/n2910 , 
        \ALUSHT/SHT/n2880 , \ALUSHT/SHT/n2749 , \ALUSHT/SHT/n2373 , 
        \ALUSHT/SHT/n2562 , \ALUSHT/SHT/n2479 , \ALUSHT/SHT/n2810 , 
        \ALUSHT/SHT/n2752 , \ALUSHT/SHT/n2462 , \ALUSHT/SHT/n2980 , 
        \ALUSHT/SHT/n2965 , \ALUSHT/SHT/n2445 , \ALUSHT/SHT/n3110 , 
        \ALUSHT/SHT/n2837 , \ALUSHT/SHT/n3080 , \ALUSHT/SHT/n2368 , 
        \ALUSHT/SHT/n2321 , \ALUSHT/SHT/n2649 , \ALUSHT/SHT/n2579 , 
        \ALUSHT/SHT/n2790 , \ALUSHT/SHT/n3065 , \ALUSHT/SHT/n2600 , 
        \ALUSHT/SHT/n2942 , \ALUSHT/SHT/n2530 , \ALUSHT/SHT/n2306 , 
        \ALUSHT/SHT/n2517 , \ALUSHT/SHT/n2627 , \ALUSHT/SHT/n2487 , 
        \ALUSHT/SHT/n3042 , \ALUSHT/SHT/n2859 , \ALUSHT/SHT/n2919 , 
        \ALUSHT/SHT/n2505 , \ALUSHT/SHT/n2439 , \ALUSHT/SHT/n2699 , 
        \ALUSHT/SHT/n2709 , \ALUSHT/SHT/n2612 , \ALUSHT/SHT/n3077 , 
        \ALUSHT/SHT/n2495 , \ALUSHT/SHT/n2314 , \ALUSHT/SHT/n2333 , 
        \ALUSHT/SHT/n2522 , \ALUSHT/SHT/n2782 , \ALUSHT/SHT/n2950 , 
        \ALUSHT/SHT/n2635 , \ALUSHT/SHT/n2977 , \ALUSHT/SHT/n3050 , 
        \ALUSHT/SHT/n2889 , \ALUSHT/SHT/n3019 , \ALUSHT/SHT/n2457 , 
        \ALUSHT/SHT/n2740 , \ALUSHT/SHT/n2470 , \ALUSHT/SHT/n2802 , 
        \ALUSHT/SHT/n2992 , \ALUSHT/SHT/n2767 , \ALUSHT/SHT/n3092 , 
        \ALUSHT/SHT/n3102 , \ALUSHT/SHT/n2825 , \ALUSHT/SHT/n2925 , 
        \ALUSHT/SHT/n2819 , \ALUSHT/SHT/n2989 , \ALUSHT/SHT/n3089 , 
        \ALUSHT/SHT/n2346 , \ALUSHT/SHT/n2557 , \ALUSHT/SHT/n2532 , 
        \ALUSHT/SHT/n2667 , \ALUSHT/SHT/n2570 , \ALUSHT/SHT/n2640 , 
        \ALUSHT/SHT/n3002 , \ALUSHT/SHT/n3025 , \ALUSHT/SHT/n2539 , 
        \ALUSHT/SHT/n2902 , \ALUSHT/SHT/n2361 , \ALUSHT/SHT/n2892 , 
        \ALUSHT/SHT/n2735 , \ALUSHT/SHT/n2328 , \ALUSHT/SHT/n2799 , 
        \ALUSHT/SHT/n2609 , \ALUSHT/SHT/n2682 , \ALUSHT/SHT/n2877 , 
        \ALUSHT/SHT/n2384 , \ALUSHT/SHT/n2405 , \ALUSHT/SHT/n2595 , 
        \ALUSHT/SHT/n2422 , \ALUSHT/SHT/n2850 , \ALUSHT/SHT/n2689 , 
        \ALUSHT/SHT/n2712 , \ALUSHT/SHT/n2719 , \ALUSHT/SHT/n2323 , 
        \ALUSHT/SHT/n2967 , \ALUSHT/SHT/n2304 , \ALUSHT/SHT/n2429 , 
        \ALUSHT/SHT/n2515 , \ALUSHT/SHT/n2485 , \ALUSHT/SHT/n2792 , 
        \ALUSHT/SHT/n2625 , \ALUSHT/SHT/n3040 , \ALUSHT/SHT/n2602 , 
        \ALUSHT/SHT/n3067 , \ALUSHT/SHT/n2940 , \ALUSHT/SHT/n3009 , 
        \ALUSHT/SHT/n2982 , \ALUSHT/SHT/n2460 , \ALUSHT/SHT/n2447 , 
        \ALUSHT/SHT/n2899 , \ALUSHT/SHT/n2777 , \ALUSHT/SHT/n2909 , 
        \ALUSHT/SHT/n3082 , \ALUSHT/SHT/n2835 , \ALUSHT/SHT/n2812 , 
        \ALUSHT/SHT/n2750 , \ALUSHT/SHT/n2809 , \ALUSHT/SHT/n2999 , 
        \ALUSHT/SHT/n3109 , \ALUSHT/SHT/n3099 , \ALUSHT/SHT/n2927 , 
        \ALUSHT/SHT/n2386 , \ALUSHT/SHT/n2529 , \ALUSHT/SHT/n2650 , 
        \ALUSHT/SHT/n3035 , \ALUSHT/SHT/n2882 , \ALUSHT/SHT/n2371 , 
        \ALUSHT/SHT/n2560 , \ALUSHT/SHT/n2547 , \ALUSHT/SHT/n2912 , 
        \ALUSHT/SHT/n2356 , \ALUSHT/SHT/n2935 , \ALUSHT/SHT/n3012 , 
        \ALUSHT/SHT/n2338 , \ALUSHT/SHT/n2677 , \ALUSHT/SHT/n2737 , 
        \ALUSHT/SHT/n2692 , \ALUSHT/SHT/n2619 , \ALUSHT/SHT/n2789 , 
        \ALUSHT/SHT/n2702 , \ALUSHT/SHT/n2432 , \ALUSHT/SHT/n2840 , 
        \ALUSHT/SHT/n2852 , \ALUSHT/SHT/n2725 , \ALUSHT/SHT/n2867 , 
        \ALUSHT/SHT/n2585 , \ALUSHT/SHT/n2415 , \ALUSHT/SHT/n2394 , 
        \ALUSHT/SHT/n2420 , \ALUSHT/SHT/n2680 , \ALUSHT/SHT/n2710 , 
        \ALUSHT/SHT/n2875 , \ALUSHT/SHT/n2949 , \ALUSHT/SHT/n2407 , 
        \ALUSHT/SHT/n2597 , \ALUSHT/SHT/n3027 , \ALUSHT/SHT/n3049 , 
        \ALUSHT/SHT/n2900 , \ALUSHT/SHT/n2642 , \ALUSHT/SHT/n2890 , 
        \ALUSHT/SHT/n2363 , \ALUSHT/SHT/n2572 , \ALUSHT/SHT/n2759 , 
        \ALUSHT/SHT/n2344 , \ALUSHT/SHT/n2555 , \ALUSHT/SHT/n2665 , 
        \ALUSHT/SHT/n3000 , \ALUSHT/SHT/n2469 , \ALUSHT/SHT/n2952 , 
        \ALUSHT/SHT/n2780 , \ALUSHT/SHT/n2316 , \ALUSHT/SHT/n2975 , 
        \ALUSHT/SHT/n2378 , \ALUSHT/SHT/n2765 , \ALUSHT/SHT/n3090 , 
        \ALUSHT/SHT/n3100 , \ALUSHT/SHT/n2455 , \ALUSHT/SHT/n2827 , 
        \ALUSHT/SHT/n2472 , \ALUSHT/SHT/n2800 , \ALUSHT/SHT/n2990 , 
        \ALUSHT/SHT/n2569 , \ALUSHT/SHT/n2742 , \ALUSHT/SHT/n2659 , 
        \ALUSHT/SHT/n2497 , \ALUSHT/SHT/n2507 , \ALUSHT/SHT/n2610 , 
        \ALUSHT/SHT/n2637 , \ALUSHT/SHT/n3052 , \ALUSHT/SHT/n3075 , 
        \ALUSHT/SHT/n2331 , \ALUSHT/SHT/n2520 , \ALUSHT/SHT/n2617 , 
        \ALUSHT/SHT/n2849 , \ALUSHT/SHT/n2955 , \ALUSHT/SHT/n2336 , 
        \ALUSHT/SHT/n2527 , \ALUSHT/SHT/n3072 , \ALUSHT/SHT/n2787 , 
        \ALUSHT/SHT/n2490 , \ALUSHT/SHT/n2500 , \ALUSHT/SHT/n3055 , 
        \ALUSHT/SHT/n2630 , \ALUSHT/SHT/n2311 , \ALUSHT/SHT/n2972 , 
        \ALUSHT/SHT/n2400 , \ALUSHT/SHT/n2920 , \ALUSHT/SHT/n2807 , 
        \ALUSHT/SHT/n2745 , \ALUSHT/SHT/n2869 , \ALUSHT/SHT/n2475 , 
        \ALUSHT/SHT/n2549 , \ALUSHT/SHT/n2762 , \ALUSHT/SHT/n2452 , 
        \ALUSHT/SHT/n2997 , \ALUSHT/SHT/n2820 , \ALUSHT/SHT/n3097 , 
        \ALUSHT/SHT/n3107 , \ALUSHT/SHT/n2662 , \ALUSHT/SHT/n2358 , 
        \ALUSHT/SHT/n2679 , \ALUSHT/SHT/n2343 , \ALUSHT/SHT/n2552 , 
        \ALUSHT/SHT/n3007 , \ALUSHT/SHT/n2897 , \ALUSHT/SHT/n2364 , 
        \ALUSHT/SHT/n2575 , \ALUSHT/SHT/n2645 , \ALUSHT/SHT/n2907 , 
        \ALUSHT/SHT/n2779 , \ALUSHT/SHT/n3020 , \ALUSHT/SHT/n2449 , 
        \ALUSHT/SHT/n2590 , \ALUSHT/SHT/n2393 , \ALUSHT/SHT/n2381 , 
        \ALUSHT/SHT/n2639 , \ALUSHT/SHT/n2730 , \ALUSHT/SHT/n2872 , 
        \ALUSHT/SHT/n2318 , \ALUSHT/SHT/n2427 , \ALUSHT/SHT/n2687 , 
        \ALUSHT/SHT/n2717 , \ALUSHT/SHT/n2969 , \ALUSHT/SHT/n2855 , 
        \ALUSHT/SHT/n2499 , \ALUSHT/SHT/n3069 , \ALUSHT/SHT/n2509 , 
        \ALUSHT/SHT/n2860 , \ALUSHT/SHT/n2412 , \ALUSHT/SHT/n2435 , 
        \ALUSHT/SHT/n2847 , \ALUSHT/SHT/n2722 , \ALUSHT/SHT/n2582 , 
        \ALUSHT/SHT/n2695 , \ALUSHT/SHT/n2705 , \ALUSHT/SHT/n2829 , 
        \ALUSHT/SHT/n2915 , \ALUSHT/SHT/n2540 , \ALUSHT/SHT/n2670 , 
        \ALUSHT/SHT/n2351 , \ALUSHT/SHT/n2932 , \ALUSHT/SHT/n3015 , 
        \ALUSHT/SHT/n2885 , \ALUSHT/SHT/n2376 , \ALUSHT/SHT/n2567 , 
        \ALUSHT/SHT/n2657 , \ALUSHT/SHT/n3029 , \ALUSHT/SHT/n3032 , 
        \ALUSHT/SHT/n2388 , \ALUSHT/SHT/n2929 , \ALUSHT/SHT/n2409 , 
        \ALUSHT/SHT/n2440 , \ALUSHT/SHT/n2757 , \ALUSHT/SHT/n2467 , 
        \ALUSHT/SHT/n2815 , \ALUSHT/SHT/n2985 , \ALUSHT/SHT/n2832 , 
        \ALUSHT/SHT/n2739 , \ALUSHT/SHT/n2770 , \ALUSHT/SHT/n3085 , 
        \ALUSHT/SHT/n2401 , \ALUSHT/SHT/n2303 , \ALUSHT/SHT/n2795 , 
        \ALUSHT/SHT/n2324 , \ALUSHT/SHT/n2947 , \ALUSHT/SHT/n2599 , 
        \ALUSHT/SHT/n2535 , \ALUSHT/SHT/n2605 , \ALUSHT/SHT/n3060 , 
        \ALUSHT/SHT/n2960 , \ALUSHT/SHT/n2622 , \ALUSHT/SHT/n3047 , 
        \ALUSHT/SHT/n2482 , \ALUSHT/SHT/n2380 , \ALUSHT/SHT/n2512 , 
        \ALUSHT/SHT/n2631 , \ALUSHT/SHT/n2526 , \ALUSHT/SHT/n2548 , 
        \ALUSHT/SHT/n2574 , \ALUSHT/SHT/n2921 , \ALUSHT/SHT/n2873 , 
        \ALUSHT/SHT/n2591 , \ALUSHT/SHT/n2854 , \ALUSHT/SHT/n2686 , 
        \ALUSHT/SHT/n2731 , \ALUSHT/SHT/n2426 , \ALUSHT/SHT/n2716 , 
        \ALUSHT/SHT/n2342 , \ALUSHT/SHT/n2663 , \ALUSHT/SHT/n2968 , 
        \ALUSHT/SHT/n3006 , \ALUSHT/SHT/n3068 , \ALUSHT/SHT/n2553 , 
        \ALUSHT/SHT/n2778 , \ALUSHT/SHT/n2644 , \ALUSHT/SHT/n2896 , 
        \ALUSHT/SHT/n2365 , \ALUSHT/SHT/n2906 , \ALUSHT/SHT/n3021 , 
        \ALUSHT/SHT/n2744 , \ALUSHT/SHT/n2448 , \ALUSHT/SHT/n2763 , 
        \ALUSHT/SHT/n2806 , \ALUSHT/SHT/n2474 , \ALUSHT/SHT/n2996 , 
        \ALUSHT/SHT/n2453 , \ALUSHT/SHT/n2821 , \ALUSHT/SHT/n3096 , 
        \ALUSHT/SHT/n3106 , \ALUSHT/SHT/n2359 , \ALUSHT/SHT/n2678 , 
        \ALUSHT/SHT/n2954 , \ALUSHT/SHT/n2337 , \ALUSHT/SHT/n2616 , 
        \ALUSHT/SHT/n2786 , \ALUSHT/SHT/n3073 , \ALUSHT/SHT/n2491 , 
        \ALUSHT/SHT/n2310 , \ALUSHT/SHT/n3054 , \ALUSHT/SHT/n2973 , 
        \ALUSHT/SHT/n2501 , \ALUSHT/SHT/n2389 , \ALUSHT/SHT/n2738 , 
        \ALUSHT/SHT/n2868 , \ALUSHT/SHT/n2598 , \ALUSHT/SHT/n2928 , 
        \ALUSHT/SHT/n3046 , \ALUSHT/SHT/n2946 , \ALUSHT/SHT/n2408 , 
        \ALUSHT/SHT/n2794 , \ALUSHT/SHT/n2325 , \ALUSHT/SHT/n2534 , 
        \ALUSHT/SHT/n2604 , \ALUSHT/SHT/n2623 , \ALUSHT/SHT/n3061 , 
        \ALUSHT/SHT/n2302 , \ALUSHT/SHT/n2513 , \ALUSHT/SHT/n2961 , 
        \ALUSHT/SHT/n2483 , \ALUSHT/SHT/n3028 , \ALUSHT/SHT/n2441 , 
        \ALUSHT/SHT/n2814 , \ALUSHT/SHT/n2756 , \ALUSHT/SHT/n2466 , 
        \ALUSHT/SHT/n2984 , \ALUSHT/SHT/n2833 , \ALUSHT/SHT/n3084 , 
        \ALUSHT/SHT/n2828 , \ALUSHT/SHT/n2771 , \ALUSHT/SHT/n2392 , 
        \ALUSHT/SHT/n2541 , \ALUSHT/SHT/n2671 , \ALUSHT/SHT/n3014 , 
        \ALUSHT/SHT/n2933 , \ALUSHT/SHT/n2566 , \ALUSHT/SHT/n2884 , 
        \ALUSHT/SHT/n2350 , \ALUSHT/SHT/n2377 , \ALUSHT/SHT/n2914 , 
        \ALUSHT/SHT/n2498 , \ALUSHT/SHT/n2656 , \ALUSHT/SHT/n3033 , 
        \ALUSHT/SHT/n2319 , \ALUSHT/SHT/n2508 , \ALUSHT/SHT/n2861 , 
        \ALUSHT/SHT/n2638 , \ALUSHT/SHT/n2583 , \ALUSHT/SHT/n2395 , 
        \ALUSHT/SHT/n2618 , \ALUSHT/SHT/n2434 , \ALUSHT/SHT/n2694 , 
        \ALUSHT/SHT/n2723 , \ALUSHT/SHT/n2413 , \ALUSHT/SHT/n2704 , 
        \ALUSHT/SHT/n2846 , \ALUSHT/SHT/n2528 , \ALUSHT/SHT/n2339 , 
        \ALUSHT/SHT/n2788 , \ALUSHT/SHT/n2724 , \ALUSHT/SHT/n2693 , 
        \ALUSHT/SHT/n2433 , \ALUSHT/SHT/n2841 , \ALUSHT/SHT/n2703 , 
        \ALUSHT/SHT/n2414 , \ALUSHT/SHT/n3108 , \ALUSHT/SHT/n2584 , 
        \ALUSHT/SHT/n2866 , \ALUSHT/SHT/n2808 , \ALUSHT/SHT/n2998 , 
        \ALUSHT/SHT/n3098 , \ALUSHT/SHT/n2651 , \ALUSHT/SHT/n2883 , 
        \ALUSHT/SHT/n2370 , \ALUSHT/SHT/n2561 , \ALUSHT/SHT/n3034 , 
        \ALUSHT/SHT/n2913 , \ALUSHT/SHT/n2546 , \ALUSHT/SHT/n2357 , 
        \ALUSHT/SHT/n2676 , \ALUSHT/SHT/n2934 , \ALUSHT/SHT/n3008 , 
        \ALUSHT/SHT/n3013 , \ALUSHT/SHT/n2506 , \ALUSHT/SHT/n2776 , 
        \ALUSHT/SHT/n2908 , \ALUSHT/SHT/n2898 , \ALUSHT/SHT/n2983 , 
        \ALUSHT/SHT/n2446 , \ALUSHT/SHT/n3083 , \ALUSHT/SHT/n2461 , 
        \ALUSHT/SHT/n2834 , \ALUSHT/SHT/n2966 , \ALUSHT/SHT/n2751 , 
        \ALUSHT/SHT/n2813 , \ALUSHT/SHT/n2305 , \ALUSHT/SHT/n2428 , 
        \ALUSHT/SHT/n2688 , \ALUSHT/SHT/n2718 , \ALUSHT/SHT/n2484 , 
        \ALUSHT/SHT/n2514 , \ALUSHT/SHT/n2974 , \ALUSHT/SHT/n2322 , 
        \ALUSHT/SHT/n2793 , \ALUSHT/SHT/n2603 , \ALUSHT/SHT/n2624 , 
        \ALUSHT/SHT/n3041 , \ALUSHT/SHT/n3066 , \ALUSHT/SHT/n2533 , 
        \ALUSHT/SHT/n2941 , \ALUSHT/SHT/n2953 , \ALUSHT/SHT/n2781 , 
        \ALUSHT/SHT/n2317 , \ALUSHT/SHT/n2496 , \ALUSHT/SHT/n2636 , 
        \ALUSHT/SHT/n3053 , \ALUSHT/SHT/n3074 , \ALUSHT/SHT/n2611 , 
        \ALUSHT/SHT/n2330 , \ALUSHT/SHT/n2521 , \ALUSHT/SHT/n2926 , 
        \ALUSHT/SHT/n3026 , \ALUSHT/SHT/n2643 , \ALUSHT/SHT/n2743 , 
        \ALUSHT/SHT/n2848 , \ALUSHT/SHT/n2801 , \ALUSHT/SHT/n2454 , 
        \ALUSHT/SHT/n2764 , \ALUSHT/SHT/n2826 , \ALUSHT/SHT/n3091 , 
        \ALUSHT/SHT/n3101 , \ALUSHT/SHT/n2473 , \ALUSHT/SHT/n2991 , 
        \ALUSHT/SHT/n2379 , \ALUSHT/SHT/n2568 , \ALUSHT/SHT/n2658 , 
        \ALUSHT/SHT/n2891 , \ALUSHT/SHT/n2901 , \ALUSHT/SHT/n2362 , 
        \ALUSHT/SHT/n2573 , \ALUSHT/SHT/n2664 , \ALUSHT/SHT/n2345 , 
        \ALUSHT/SHT/n2554 , \ALUSHT/SHT/n2853 , \ALUSHT/SHT/n2758 , 
        \ALUSHT/SHT/n3001 , \ALUSHT/SHT/n2468 , \ALUSHT/SHT/n2736 , 
        \ALUSHT/SHT/n2681 , \ALUSHT/SHT/n2421 , \ALUSHT/SHT/n2711 , 
        \ALUSHT/SHT/n2406 , \ALUSHT/SHT/n2596 , \ALUSHT/SHT/n2874 , 
        \ALUSHT/SHT/n2948 , \ALUSHT/SHT/n3048 , \REG_2/ph8dec_2/n20 , 
        \REG_2/ph8dec_2/n21 , \CODEQ/phque34_1/n753 , \CODEQ/phque34_1/n758 , 
        \CODEQ/phque34_1/n764 , \CODEQ/phque34_1/stream3[36] , 
        \CODEQ/phque34_1/n756 , \CODEQ/phque34_1/stream3[39] , 
        \CODEQ/phque34_1/n761 , \CODEQ/phque34_1/n754 , \CODEQ/phque34_1/n755 , 
        \CODEQ/phque34_1/n759 , \CODEQ/phque34_1/n757 , \CODEQ/phque34_1/n763 , 
        \CODEQ/phque34_1/n762 , \CODEQ/phque34_1/n765 , \CODEQ/phque34_1/n760 , 
        \CODEQ/phque34_1/stream3[35] , \CODEQ/phque34_1/stream3[38] , 
        \CODEQ/phque34_1/n766 , \CODEQ/phque34_1/stream3[37] , 
        \MCD/rd_wt_1/n4441 , \MCD/rd_wt_1/n4466 , \MCD/rd_wt_1/n4426 , 
        \MCD/rd_wt_1/n4434 , \MCD/rd_wt_1/n4448 , \MCD/rd_wt_1/n4453 , 
        \MCD/rd_wt_1/n4454 , \MCD/rd_wt_1/n4419 , \MCD/rd_wt_1/n4420 , 
        \MCD/rd_wt_1/n4421 , \MCD/rd_wt_1/n4428 , \MCD/rd_wt_1/n4433 , 
        \MCD/rd_wt_1/n4468 , \MCD/rd_wt_1/n4446 , \MCD/rd_wt_1/n4461 , 
        \MCD/rd_wt_1/ciff , \MCD/rd_wt_1/n4429 , \MCD/rd_wt_1/n4447 , 
        \MCD/rd_wt_1/n4455 , \MCD/rd_wt_1/n4460 , \MCD/rd_wt_1/n4432 , 
        \MCD/rd_wt_1/n4435 , \MCD/rd_wt_1/n4440 , \MCD/rd_wt_1/n4467 , 
        \MCD/rd_wt_1/n4425 , \MCD/rd_wt_1/bacc , \MCD/rd_wt_1/n4452 , 
        \MCD/rd_wt_1/n4427 , \MCD/rd_wt_1/n4437 , \MCD/rd_wt_1/n4442 , 
        \MCD/rd_wt_1/n4449 , \MCD/rd_wt_1/n4465 , \MCD/rd_wt_1/n4459 , 
        \MCD/rd_wt_1/n4422 , \MCD/rd_wt_1/n4439 , \MCD/rd_wt_1/n4450 , 
        \MCD/rd_wt_1/n4457 , \MCD/rd_wt_1/n4430 , \MCD/rd_wt_1/n4423 , 
        \MCD/rd_wt_1/n4445 , \MCD/rd_wt_1/n4462 , \MCD/rd_wt_1/n4438 , 
        \MCD/rd_wt_1/n4444 , \MCD/rd_wt_1/n4456 , \MCD/rd_wt_1/n4463 , 
        \MCD/rd_wt_1/n4431 , \MCD/rd_wt_1/n4418 , \MCD/rd_wt_1/n4436 , 
        \MCD/rd_wt_1/n4458 , \MCD/rd_wt_1/n4443 , \MCD/rd_wt_1/n4451 , 
        \MCD/rd_wt_1/n4464 , \MCD/rd_wt_1/n4424 , \MAIN/STM/exec_eoc , 
        \MAIN/STM/exe_1st_r , \MAIN/STM/seq_doing , \MAIN/STM/exec_eoc1 , 
        \MAIN/STM/exec_end3 , \MAIN/STM/seq_end , \MAIN/STM/n3366 , 
        \MAIN/STM/exe_1st , \MAIN/STM/exe_2nd , \MAIN/STM/exe_err2 , 
        \MAIN/STM/exe_1st_w , \MAIN/STM/exe_2nd_w , \MAIN/STM/sa_start3 , 
        \MAIN/STM/exe_err3 , \MAIN/STM/exec_end2 , \MAIN/STM/sa_start2 , 
        \MAIN/STM/srgfilewren_h , \MAIN/STM/exec_eoc2 , \MAIN/STM/n3365 , 
        \MAIN/STM/bnolth , \MAIN/STM/exestage_err , \MAIN/STM/execute_err , 
        \MAIN/STM/exec_end1 , \MAIN/STM/n3364 , \MAIN/STM/exec_eoc3 , 
        \MAIN/SW/nst[0] , \MAIN/SW/wst[0] , \MAIN/SW/n3322 , \MAIN/SW/n3323 , 
        \CODEQ/phque12_1/n767 , \CODEQ/phque12_1/n771 , 
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 , \CODEQ/phque12_1/queue2[22] , 
        \CODEQ/phque12_1/queue2[18] , \CODEQ/phque12_1/queue2[11] , 
        \CODEQ/phque12_1/queue2[26] , \CODEQ/phque12_1/queue2[6] , 
        \CODEQ/phque12_1/queue1[5] , \CODEQ/phque12_1/queue2[15] , 
        \CODEQ/phque12_1/queue1[56] , \CODEQ/phque12_1/queue1[8] , 
        \CODEQ/phque12_1/queue2[2] , \CODEQ/phque12_1/queue1[1] , 
        \CODEQ/phque12_1/queue2[36] , \CODEQ/phque12_1/queue2[0] , 
        \CODEQ/phque12_1/queue1[3] , \CODEQ/phque12_1/queue2[9] , 
        \CODEQ/phque12_1/queue2[24] , \CODEQ/phque12_1/queue2[17] , 
        \CODEQ/phque12_1/queue2[4] , \CODEQ/phque12_1/queue1[7] , 
        \CODEQ/phque12_1/n770 , \CODEQ/phque12_1/queue2[39] , 
        \CODEQ/phque12_1/queue2[30] , \CODEQ/phque12_1/queue2[29] , 
        \CODEQ/phque12_1/queue1[40] , \CODEQ/phque12_1/queue1[49] , 
        \CODEQ/phque12_1/queue2[20] , \CODEQ/phque12_1/queue2[13] , 
        \CODEQ/phque12_1/queue1[35] , \CODEQ/phque12_1/queue2[55] , 
        \CODEQ/phque12_1/queue1[25] , \CODEQ/phque12_1/queue1[16] , 
        \CODEQ/phque12_1/queue1[31] , \CODEQ/phque12_1/queue1[28] , 
        \CODEQ/phque12_1/queue2[48] , \CODEQ/phque12_1/queue1[38] , 
        \CODEQ/phque12_1/queue1[12] , \CODEQ/phque12_1/queue1[21] , 
        \CODEQ/phque12_1/queue1[23] , \CODEQ/phque12_1/queue1[10] , 
        \CODEQ/phque12_1/queue1[19] , \CODEQ/phque12_1/queue1[27] , 
        \CODEQ/phque12_1/queue1[14] , \CODEQ/phque12_1/queue2[56] , 
        \CODEQ/phque12_1/queue1[37] , \CODEQ/phque12_1/queue1[26] , 
        \CODEQ/phque12_1/queue1[15] , \CODEQ/phque12_1/n769 , 
        \CODEQ/phque12_1/queue1[36] , \CODEQ/phque12_1/queue1[22] , 
        \CODEQ/phque12_1/queue1[11] , \CODEQ/phque12_1/queue1[18] , 
        \CODEQ/phque12_1/queue2[40] , \CODEQ/phque12_1/queue2[49] , 
        \CODEQ/phque12_1/queue1[39] , \CODEQ/phque12_1/queue1[30] , 
        \CODEQ/phque12_1/queue1[29] , \CODEQ/phque12_1/queue1[20] , 
        \CODEQ/phque12_1/queue1[13] , \CODEQ/phque12_1/n768 , 
        \CODEQ/phque12_1/queue1[24] , \CODEQ/phque12_1/queue1[17] , 
        \CODEQ/phque12_1/queue2[5] , \CODEQ/phque12_1/queue1[6] , 
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 , \CODEQ/phque12_1/queue2[38] , 
        \CODEQ/phque12_1/queue2[31] , \CODEQ/phque12_1/queue2[28] , 
        \CODEQ/phque12_1/queue2[21] , \CODEQ/phque12_1/queue2[12] , 
        \CODEQ/phque12_1/queue1[48] , \CODEQ/phque12_1/queue2[35] , 
        \CODEQ/phque12_1/queue2[1] , \CODEQ/phque12_1/queue1[2] , 
        \CODEQ/phque12_1/queue2[8] , \CODEQ/phque12_1/queue2[27] , 
        \CODEQ/phque12_1/queue2[25] , \CODEQ/phque12_1/queue1[55] , 
        \CODEQ/phque12_1/queue2[16] , \CODEQ/phque12_1/queue2[14] , 
        \CODEQ/phque12_1/queue1[9] , \CODEQ/phque12_1/queue2[3] , 
        \CODEQ/phque12_1/queue1[0] , \CODEQ/phque12_1/queue2[37] , 
        \CODEQ/phque12_1/queue2[23] , \CODEQ/phque12_1/queue2[19] , 
        \CODEQ/phque12_1/queue2[10] , \CODEQ/phque12_1/queue2[7] , 
        \CODEQ/phque12_1/queue1[4] , \SADR/SELSEG/n9104 , \SADR/SELSEG/n9087 , 
        \SADR/SELSEG/n8945 , \SADR/SELSEG/n8962 , \SADR/SELSEG/n9045 , 
        \SADR/SELSEG/n9062 , \SADR/SELSEG/n9092 , \SADR/SELSEG/n9117 , 
        \SADR/SELSEG/n9105 , \SADR/SELSEG/n8930 , \SADR/SELSEG/n8987 , 
        \SADR/SELSEG/n9030 , \SADR/SELSEG/n8979 , \SADR/SELSEG/n9017 , 
        \SADR/SELSEG/n9079 , \SADR/SELSEG/n9005 , \SADR/SELSEG/n9022 , 
        \SADR/SELSEG/n9095 , \SADR/SELSEG/n8939 , \SADR/SELSEG/n8995 , 
        \SADR/SELSEG/n8950 , \SADR/SELSEG/n8957 , \SADR/SELSEG/n8970 , 
        \SADR/SELSEG/n9039 , \SADR/SELSEG/n9057 , \SADR/SELSEG/n9070 , 
        \SADR/SELSEG/n8977 , \SADR/SELSEG/n9050 , \SADR/SELSEG/n9077 , 
        \SADR/SELSEG/n8992 , \SADR/SELSEG/n9102 , \SADR/SELSEG/n9089 , 
        \SADR/SELSEG/n9002 , \SADR/SELSEG/n9019 , \SADR/SELSEG/n9025 , 
        \SADR/SELSEG/n9076 , \SADR/SELSEG/n9110 , \SADR/SELSEG/n8937 , 
        \SADR/SELSEG/n8959 , \SADR/SELSEG/n8989 , \SADR/SELSEG/n9059 , 
        \SADR/SELSEG/n9010 , \SADR/SELSEG/n8980 , \SADR/SELSEG/n9037 , 
        \SADR/SELSEG/n9080 , \SADR/SELSEG/n8942 , \SADR/SELSEG/n8965 , 
        \SADR/SELSEG/n9042 , \SADR/SELSEG/n9065 , \SADR/SELSEG/n8988 , 
        \SADR/SELSEG/n9003 , \SADR/SELSEG/n9024 , \SADR/SELSEG/n9088 , 
        \SADR/SELSEG/n9118 , \SADR/SELSEG/n8951 , \SADR/SELSEG/n8993 , 
        \SADR/SELSEG/n9093 , \SADR/SELSEG/n9103 , \SADR/SELSEG/n9018 , 
        \SADR/SELSEG/n9094 , \SADR/SELSEG/n9078 , \SADR/SELSEG/n9111 , 
        \SADR/SELSEG/n8976 , \SADR/SELSEG/n9051 , \SADR/SELSEG/n8943 , 
        \SADR/SELSEG/n8964 , \SADR/SELSEG/n9064 , \SADR/SELSEG/n9043 , 
        \SADR/SELSEG/n8981 , \SADR/SELSEG/n9081 , \SADR/SELSEG/n8936 , 
        \SADR/SELSEG/n9011 , \SADR/SELSEG/n8958 , \SADR/SELSEG/n9036 , 
        \SADR/SELSEG/n9058 , \SADR/SELSEG/n9086 , \SADR/SELSEG/n9116 , 
        \SADR/SELSEG/n8931 , \SADR/SELSEG/n8978 , \SADR/SELSEG/n9031 , 
        \SADR/SELSEG/n9016 , \SADR/SELSEG/n8986 , \SADR/SELSEG/n8944 , 
        \SADR/SELSEG/n8963 , \SADR/SELSEG/n9044 , \SADR/SELSEG/n9063 , 
        \SADR/SELSEG/n8956 , \SADR/SELSEG/n8971 , \SADR/SELSEG/n9056 , 
        \SADR/SELSEG/n9071 , \SADR/SELSEG/n9084 , \SADR/SELSEG/n9114 , 
        \SADR/SELSEG/n8938 , \SADR/SELSEG/n8994 , \SADR/SELSEG/n9004 , 
        \SADR/SELSEG/n9023 , \SADR/SELSEG/n9038 , \SADR/SELSEG/n8946 , 
        \SADR/SELSEG/n9061 , \SADR/SELSEG/n8961 , \SADR/SELSEG/n8984 , 
        \SADR/SELSEG/n9046 , \SADR/SELSEG/n9109 , \SADR/SELSEG/n9112 , 
        \SADR/SELSEG/n9090 , \SADR/SELSEG/n9091 , \SADR/SELSEG/n9106 , 
        \SADR/SELSEG/n9096 , \SADR/SELSEG/n8933 , \SADR/SELSEG/n9028 , 
        \SADR/SELSEG/n9014 , \SADR/SELSEG/n9033 , \SADR/SELSEG/n8968 , 
        \SADR/SELSEG/n9006 , \SADR/SELSEG/n9068 , \SADR/SELSEG/n9021 , 
        \SADR/SELSEG/n8996 , \SADR/SELSEG/n9101 , \SADR/SELSEG/n8954 , 
        \SADR/SELSEG/n9073 , \SADR/SELSEG/n8973 , \SADR/SELSEG/n9054 , 
        \SADR/SELSEG/n8953 , \SADR/SELSEG/n8974 , \SADR/SELSEG/n9053 , 
        \SADR/SELSEG/n9074 , \SADR/SELSEG/n8948 , \SADR/SELSEG/n8991 , 
        \SADR/SELSEG/n9001 , \SADR/SELSEG/n9026 , \SADR/SELSEG/n9048 , 
        \SADR/SELSEG/n8934 , \SADR/SELSEG/n9034 , \SADR/SELSEG/n9013 , 
        \SADR/SELSEG/n8941 , \SADR/SELSEG/n8966 , \SADR/SELSEG/n8983 , 
        \SADR/SELSEG/n8998 , \SADR/SELSEG/n9083 , \SADR/SELSEG/n9098 , 
        \SADR/SELSEG/n9108 , \SADR/SELSEG/n9113 , \SADR/SELSEG/n9008 , 
        \SADR/SELSEG/n9041 , \SADR/SELSEG/n9066 , \SADR/SELSEG/n8949 , 
        \SADR/SELSEG/n9000 , \SADR/SELSEG/n9027 , \SADR/SELSEG/n9049 , 
        \SADR/SELSEG/n9100 , \SADR/SELSEG/n8940 , \SADR/SELSEG/n8952 , 
        \SADR/SELSEG/n8975 , \SADR/SELSEG/n8990 , \SADR/SELSEG/n9052 , 
        \SADR/SELSEG/n8967 , \SADR/SELSEG/n9040 , \SADR/SELSEG/n9075 , 
        \SADR/SELSEG/n9067 , \SADR/SELSEG/n9082 , \SADR/SELSEG/n8935 , 
        \SADR/SELSEG/n8982 , \SADR/SELSEG/n9009 , \SADR/SELSEG/n9012 , 
        \SADR/SELSEG/n9035 , \SADR/SELSEG/n8999 , \SADR/SELSEG/n9099 , 
        \SADR/SELSEG/n9107 , \SADR/SELSEG/n9085 , \SADR/SELSEG/n8932 , 
        \SADR/SELSEG/n8985 , \SADR/SELSEG/n9015 , \SADR/SELSEG/n9032 , 
        \SADR/SELSEG/n9115 , \SADR/SELSEG/n8929 , \SADR/SELSEG/n9029 , 
        \SADR/SELSEG/n8947 , \SADR/SELSEG/n9060 , \SADR/SELSEG/n8955 , 
        \SADR/SELSEG/n8960 , \SADR/SELSEG/n9047 , \SADR/SELSEG/n9072 , 
        \SADR/SELSEG/n8972 , \SADR/SELSEG/n8997 , \SADR/SELSEG/n9055 , 
        \SADR/SELSEG/n9097 , \SADR/SELSEG/n8969 , \SADR/SELSEG/n9007 , 
        \SADR/SELSEG/n9020 , \SADR/SELSEG/n9069 , 
        \REGF/pbmemcnt1/add_53/carry[4] , \REGF/pbmemcnt1/add_53/carry[9] , 
        \REGF/pbmemcnt1/add_53/carry[2] , \REGF/pbmemcnt1/add_53/carry[6] , 
        \REGF/pbmemcnt1/add_53/carry[11] , \REGF/pbmemcnt1/add_53/carry[10] , 
        \REGF/pbmemcnt1/add_53/carry[3] , \REGF/pbmemcnt1/add_53/carry[7] , 
        \REGF/pbmemcnt1/add_53/carry[8] , \REGF/pbmemcnt1/add_53/carry[5] , 
        \REGF/pbmemcnt1/sub_48/carry[4] , \REGF/pbmemcnt1/sub_48/carry[2] , 
        \REGF/pbmemcnt1/sub_48/carry[6] , \REGF/pbmemcnt1/sub_48/carry[7] , 
        \REGF/pbmemcnt1/sub_48/carry[3] , \REGF/pbmemcnt1/sub_48/carry[5] , 
        \REG_2/SATIME/add_187/carry[4] , \REG_2/SATIME/add_187/carry[9] , 
        \REG_2/SATIME/add_187/carry[2] , \REG_2/SATIME/add_187/carry[6] , 
        \REG_2/SATIME/add_187/carry[20] , \REG_2/SATIME/add_187/carry[13] , 
        \REG_2/SATIME/add_187/carry[17] , \REG_2/SATIME/add_187/carry[15] , 
        \REG_2/SATIME/add_187/carry[18] , \REG_2/SATIME/add_187/carry[11] , 
        \REG_2/SATIME/add_187/carry[19] , \REG_2/SATIME/add_187/carry[10] , 
        \REG_2/SATIME/add_187/carry[14] , \REG_2/SATIME/add_187/carry[16] , 
        \REG_2/SATIME/add_187/carry[12] , \REG_2/SATIME/add_187/carry[3] , 
        \REG_2/SATIME/add_187/carry[7] , \REG_2/SATIME/add_187/carry[8] , 
        \REG_2/SATIME/add_187/carry[5] , \SAEXE/RFIO/phcont4_1/ncnt[1] , 
        \SAEXE/RFIO/phcont4_1/count[0] , \SAEXE/RFIO/phcont4_1/count52[1] , 
        \SAEXE/RFIO/phcont4_1/n_42 , \SAEXE/RFIO/phcont4_1/n83 , 
        \SAEXE/RFIO/phcont4_1/ncnt[0] , \SAEXE/RFIO/phcont4_1/n84 , 
        \SAEXE/RFIO/phcont4_1/count[1] , \SAEXE/RFIO/phcont4_1/count52[0] , 
        \SAEXE/RFIO/phcont4_1/n86 , \SAEXE/RFIO/phcont4_1/n87 , 
        \SAEXE/RFIO/RIN1/nfst[2] , \SAEXE/RFIO/RIN1/n175 , 
        \SAEXE/RFIO/RIN1/n167 , \SAEXE/RFIO/RIN1/n168 , \SAEXE/RFIO/RIN1/n169 , 
        \SAEXE/RFIO/RIN1/nfst[0] , \SAEXE/RFIO/RIN1/n172 , 
        \SAEXE/RFIO/RIN1/n173 , \SAEXE/RFIO/RIN1/fst[1] , 
        \SAEXE/RFIO/RIN1/n174 , \SAEXE/RFIO/RIN1/n166 , 
        \SAEXE/RFIO/RIN1/fst[2] , \SAEXE/RFIO/RIN1/n176 , 
        \SAEXE/RFIO/RIN1/n170 , \SAEXE/RFIO/RIN1/n171 , 
        \SAEXE/RFIO/RIN1/nfst[1] , \SAEXE/RFIO/RIN1/n165 , 
        \SADR/MAINSADR/addidxof/gg_out[0] , \SADR/MAINSADR/addidxof/c_last , 
        \SADR/MAINSADR/addidxof/n8632 , \SADR/MAINSADR/addidxof/gg_out[2] , 
        \SADR/MAINSADR/addidxof/gp_out[3] , 
        \SADR/MAINSADR/addidxof/cin_stg[1] , 
        \SADR/MAINSADR/addidxof/gp_out[1] , 
        \SADR/MAINSADR/addidxof/cin_stg[2] , 
        \SADR/MAINSADR/addidxof/gp_out[2] , \SADR/MAINSADR/addidxof/gg_out[1] , 
        \SADR/MAINSADR/addidxof/gg_out[3] , 
        \SADR/MAINSADR/addsegoff/gg_out[0] , \SADR/MAINSADR/addsegoff/n8502 , 
        \SADR/MAINSADR/addsegoff/n8503 , \SADR/MAINSADR/addsegoff/gp_out[1] , 
        \SADR/MAINSADR/addsegoff/n8498 , \SADR/MAINSADR/addsegoff/n8501 , 
        \SADR/MAINSADR/addsegoff/n8497 , \SADR/MAINSADR/addsegoff/gg_out[1] , 
        \SADR/MAINSADR/addsegoff/n8499 , \SADR/MAINSADR/addsegoff/n8500 , 
        \SADR/MAINSADR/adrinc1/gg_out[4] , \SADR/MAINSADR/adrinc1/gg_out[2] , 
        \SADR/MAINSADR/adrinc1/gp_out[3] , \SADR/MAINSADR/adrinc1/gp_out[1] , 
        \SADR/MAINSADR/adrinc1/gp_out[0] , \SADR/MAINSADR/adrinc1/gp_out[4] , 
        \SADR/MAINSADR/adrinc1/gp_out[2] , \SADR/MAINSADR/adrinc1/gg_out[1] , 
        \SADR/MAINSADR/adrinc1/gg_out[3] , \SADR/MAINSADR/adrcmp1/ggfl[3] , 
        \SADR/MAINSADR/adrcmp1/n8405 , \SADR/MAINSADR/adrcmp1/ggfl[0] , 
        \SADR/MAINSADR/adrcmp1/n8404 , \SADR/MAINSADR/adrcmp1/geq[0] , 
        \SADR/MAINSADR/adrcmp1/ggfl[2] , \SADR/MAINSADR/adrcmp1/geq[2] , 
        \SADR/MAINSADR/adrcmp1/geq[3] , \SADR/MAINSADR/adrcmp1/geq[1] , 
        \SADR/MAINSADR/adrcmp1/n8406 , \SADR/MAINSADR/adrcmp1/ggfl[1] , 
        \SADR/MAINSADR/adrdec1/gg_out[0] , \SADR/MAINSADR/adrdec1/gg_out[4] , 
        \SADR/MAINSADR/adrdec1/gg_out[2] , \SADR/MAINSADR/adrdec1/gcarry[1] , 
        \SADR/MAINSADR/adrdec1/n8347 , \SADR/MAINSADR/adrdec1/gcarry[3] , 
        \SADR/MAINSADR/adrdec1/gcarry[2] , \SADR/MAINSADR/adrdec1/gcarry[4] , 
        \SADR/MAINSADR/adrdec1/gg_out[1] , \SADR/MAINSADR/adrdec1/gg_out[3] , 
        \SADR/MAINSADR/adrinc2/gg_out[4] , \SADR/MAINSADR/adrinc2/gg_out[2] , 
        \SADR/MAINSADR/adrinc2/gp_out[3] , \SADR/MAINSADR/adrinc2/gp_out[1] , 
        \SADR/MAINSADR/adrinc2/gp_out[0] , \SADR/MAINSADR/adrinc2/gp_out[4] , 
        \SADR/MAINSADR/adrinc2/gp_out[2] , \SADR/MAINSADR/adrinc2/gg_out[1] , 
        \SADR/MAINSADR/adrinc2/gg_out[3] , \SADR/MAINSADR/adrdec2/gg_out[0] , 
        \SADR/MAINSADR/adrdec2/gg_out[4] , \SADR/MAINSADR/adrdec2/gg_out[2] , 
        \SADR/MAINSADR/adrdec2/gcarry[1] , \SADR/MAINSADR/adrdec2/gcarry[3] , 
        \SADR/MAINSADR/adrdec2/n8299 , \SADR/MAINSADR/adrdec2/gcarry[2] , 
        \SADR/MAINSADR/adrdec2/gcarry[4] , \SADR/MAINSADR/adrdec2/gg_out[1] , 
        \SADR/MAINSADR/adrdec2/gg_out[3] , 
        \REGF/pbmemff21/pbinc19k_1/gg_out[2] , 
        \REGF/pbmemff21/pbinc19k_1/gp_out[3] , 
        \REGF/pbmemff21/pbinc19k_1/gp_out[1] , 
        \REGF/pbmemff21/pbinc19k_1/gp_out[0] , 
        \REGF/pbmemff21/pbinc19k_1/gp_out[2] , 
        \REGF/pbmemff21/pbinc19k_1/gg_out[3] , 
        \REGF/pbmemff21/pbinc19k_1/gg_out[1] , \SADR/ADDIDX/add_w_x/gg_out[0] , 
        \SADR/ADDIDX/add_w_x/c_last , \SADR/ADDIDX/add_w_x/gg_out[2] , 
        \SADR/ADDIDX/add_w_x/n10655 , \SADR/ADDIDX/add_w_x/gp_out[3] , 
        \SADR/ADDIDX/add_w_x/cin_stg[1] , \SADR/ADDIDX/add_w_x/gp_out[1] , 
        \SADR/ADDIDX/add_w_x/cin_stg[2] , \SADR/ADDIDX/add_w_x/gp_out[2] , 
        \SADR/ADDIDX/add_w_x/gg_out[1] , \SADR/ADDIDX/add_w_x/gg_out[3] , 
        \SADR/ADDIDX/add_x_z/gg_out[0] , \SADR/ADDIDX/add_x_z/c_last , 
        \SADR/ADDIDX/add_x_z/gg_out[2] , \SADR/ADDIDX/add_x_z/gp_out[3] , 
        \SADR/ADDIDX/add_x_z/cin_stg[1] , \SADR/ADDIDX/add_x_z/gp_out[1] , 
        \SADR/ADDIDX/add_x_z/cin_stg[2] , \SADR/ADDIDX/add_x_z/gp_out[2] , 
        \SADR/ADDIDX/add_x_z/n10526 , \SADR/ADDIDX/add_x_z/gg_out[1] , 
        \SADR/ADDIDX/add_x_z/gg_out[3] , \SADR/ADDIDX/add_y_z/gg_out[0] , 
        \SADR/ADDIDX/add_y_z/n10397 , \SADR/ADDIDX/add_y_z/c_last , 
        \SADR/ADDIDX/add_y_z/gg_out[2] , \SADR/ADDIDX/add_y_z/gp_out[3] , 
        \SADR/ADDIDX/add_y_z/cin_stg[1] , \SADR/ADDIDX/add_y_z/gp_out[1] , 
        \SADR/ADDIDX/add_y_z/cin_stg[2] , \SADR/ADDIDX/add_y_z/gp_out[2] , 
        \SADR/ADDIDX/add_y_z/gg_out[1] , \SADR/ADDIDX/add_y_z/gg_out[3] , 
        \SADR/ADDIDX/add_w_y/gg_out[0] , \SADR/ADDIDX/add_w_y/c_last , 
        \SADR/ADDIDX/add_w_y/gg_out[2] , \SADR/ADDIDX/add_w_y/gp_out[3] , 
        \SADR/ADDIDX/add_w_y/cin_stg[1] , \SADR/ADDIDX/add_w_y/gp_out[1] , 
        \SADR/ADDIDX/add_w_y/n10268 , \SADR/ADDIDX/add_w_y/cin_stg[2] , 
        \SADR/ADDIDX/add_w_y/gp_out[2] , \SADR/ADDIDX/add_w_y/gg_out[1] , 
        \SADR/ADDIDX/add_w_y/gg_out[3] , \SADR/ADDIDX/add_w_x_y/gg_out[0] , 
        \SADR/ADDIDX/add_w_x_y/c_last , \SADR/ADDIDX/add_w_x_y/gg_out[2] , 
        \SADR/ADDIDX/add_w_x_y/n10139 , \SADR/ADDIDX/add_w_x_y/gp_out[3] , 
        \SADR/ADDIDX/add_w_x_y/cin_stg[1] , \SADR/ADDIDX/add_w_x_y/gp_out[1] , 
        \SADR/ADDIDX/add_w_x_y/cin_stg[2] , \SADR/ADDIDX/add_w_x_y/gp_out[2] , 
        \SADR/ADDIDX/add_w_x_y/gg_out[1] , \SADR/ADDIDX/add_w_x_y/gg_out[3] , 
        \SADR/ADDIDX/add_x_y_z/gg_out[0] , \SADR/ADDIDX/add_x_y_z/c_last , 
        \SADR/ADDIDX/add_x_y_z/n10010 , \SADR/ADDIDX/add_x_y_z/gg_out[2] , 
        \SADR/ADDIDX/add_x_y_z/gp_out[3] , \SADR/ADDIDX/add_x_y_z/cin_stg[1] , 
        \SADR/ADDIDX/add_x_y_z/gp_out[1] , \SADR/ADDIDX/add_x_y_z/cin_stg[2] , 
        \SADR/ADDIDX/add_x_y_z/gp_out[2] , \SADR/ADDIDX/add_x_y_z/gg_out[1] , 
        \SADR/ADDIDX/add_x_y_z/gg_out[3] , \SADR/ADDIDX/add_w_z/gg_out[0] , 
        \SADR/ADDIDX/add_w_z/c_last , \SADR/ADDIDX/add_w_z/gg_out[2] , 
        \SADR/ADDIDX/add_w_z/n9881 , \SADR/ADDIDX/add_w_z/gp_out[3] , 
        \SADR/ADDIDX/add_w_z/cin_stg[1] , \SADR/ADDIDX/add_w_z/gp_out[1] , 
        \SADR/ADDIDX/add_w_z/cin_stg[2] , \SADR/ADDIDX/add_w_z/gp_out[2] , 
        \SADR/ADDIDX/add_w_z/gg_out[1] , \SADR/ADDIDX/add_w_z/gg_out[3] , 
        \SADR/ADDIDX/add_x_y/gg_out[0] , \SADR/ADDIDX/add_x_y/c_last , 
        \SADR/ADDIDX/add_x_y/gg_out[2] , \SADR/ADDIDX/add_x_y/gp_out[3] , 
        \SADR/ADDIDX/add_x_y/n9752 , \SADR/ADDIDX/add_x_y/cin_stg[1] , 
        \SADR/ADDIDX/add_x_y/gp_out[1] , \SADR/ADDIDX/add_x_y/cin_stg[2] , 
        \SADR/ADDIDX/add_x_y/gp_out[2] , \SADR/ADDIDX/add_x_y/gg_out[1] , 
        \SADR/ADDIDX/add_x_y/gg_out[3] , \SADR/ADDIDX/add_w_x_z/gg_out[0] , 
        \SADR/ADDIDX/add_w_x_z/c_last , \SADR/ADDIDX/add_w_x_z/gg_out[2] , 
        \SADR/ADDIDX/add_w_x_z/gp_out[3] , \SADR/ADDIDX/add_w_x_z/cin_stg[1] , 
        \SADR/ADDIDX/add_w_x_z/gp_out[1] , \SADR/ADDIDX/add_w_x_z/cin_stg[2] , 
        \SADR/ADDIDX/add_w_x_z/gp_out[2] , \SADR/ADDIDX/add_w_x_z/gg_out[1] , 
        \SADR/ADDIDX/add_w_x_z/gg_out[3] , \SADR/ADDIDX/add_w_x_z/n9623 , 
        \SADR/ADDIDX/add_w_y_z/gg_out[0] , \SADR/ADDIDX/add_w_y_z/c_last , 
        \SADR/ADDIDX/add_w_y_z/n9494 , \SADR/ADDIDX/add_w_y_z/gg_out[2] , 
        \SADR/ADDIDX/add_w_y_z/gp_out[3] , \SADR/ADDIDX/add_w_y_z/cin_stg[1] , 
        \SADR/ADDIDX/add_w_y_z/gp_out[1] , \SADR/ADDIDX/add_w_y_z/cin_stg[2] , 
        \SADR/ADDIDX/add_w_y_z/gp_out[2] , \SADR/ADDIDX/add_w_y_z/gg_out[1] , 
        \SADR/ADDIDX/add_w_y_z/gg_out[3] , \SADR/ADDIDX/add_w_x_y_z/gg_out[0] , 
        \SADR/ADDIDX/add_w_x_y_z/c_last , \SADR/ADDIDX/add_w_x_y_z/gg_out[2] , 
        \SADR/ADDIDX/add_w_x_y_z/gp_out[3] , 
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[1] , 
        \SADR/ADDIDX/add_w_x_y_z/gp_out[1] , 
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[2] , 
        \SADR/ADDIDX/add_w_x_y_z/gp_out[2] , 
        \SADR/ADDIDX/add_w_x_y_z/gg_out[1] , 
        \SADR/ADDIDX/add_w_x_y_z/gg_out[3] , \SADR/ADDIDX/add_w_x_y_z/n9365 , 
        \REGF/pbmemff41/phdec12_2/gg_out[0] , \REGF/pbmemff41/phdec12_2/n7080 , 
        \REGF/pbmemff41/phdec12_2/gcarry[1] , \REGF/pbmemff41/phdec12_2/n7081 , 
        \REGF/pbmemff41/phdec12_2/gg_out[1] , 
        \REGF/pbmemff41/phdec12_1/gg_out[0] , 
        \REGF/pbmemff41/phdec12_1/gcarry[1] , \REGF/pbmemff41/phdec12_1/n7063 , 
        \REGF/pbmemff41/phdec12_1/n7064 , \REGF/pbmemff41/phdec12_1/gg_out[1] , 
        \MAIN/ENGIN/STEP_A/cst[2] , \MAIN/ENGIN/STEP_A/n3545 , 
        \MAIN/ENGIN/STEP_A/n3562 , \MAIN/ENGIN/STEP_A/n3587 , 
        \MAIN/ENGIN/STEP_A/n3550 , \MAIN/ENGIN/STEP_A/n3579 , 
        \MAIN/ENGIN/STEP_A/n3557 , \MAIN/ENGIN/STEP_A/n3570 , 
        \MAIN/ENGIN/STEP_A/n3577 , \MAIN/ENGIN/STEP_A/cst[0] , 
        \MAIN/ENGIN/STEP_A/n3589 , \MAIN/ENGIN/STEP_A/tmp2[0] , 
        \MAIN/ENGIN/STEP_A/n3559 , \MAIN/ENGIN/STEP_A/n3565 , 
        \MAIN/ENGIN/STEP_A/n3580 , \MAIN/ENGIN/STEP_A/sw_stage , 
        \MAIN/ENGIN/STEP_A/n3551 , \MAIN/ENGIN/STEP_A/n3588 , 
        \MAIN/ENGIN/STEP_A/nst[3] , \MAIN/ENGIN/STEP_A/exec_stage278 , 
        \MAIN/ENGIN/STEP_A/n3576 , \MAIN/ENGIN/STEP_A/n3564 , 
        \MAIN/ENGIN/STEP_A/n3581 , \MAIN/ENGIN/STEP_A/n3558 , 
        \MAIN/ENGIN/STEP_A/n3578 , \MAIN/ENGIN/STEP_A/n3586 , 
        \MAIN/ENGIN/STEP_A/cst[3] , \MAIN/ENGIN/STEP_A/cst[1] , 
        \MAIN/ENGIN/STEP_A/n3544 , \MAIN/ENGIN/STEP_A/n3546 , 
        \MAIN/ENGIN/STEP_A/n3556 , \MAIN/ENGIN/STEP_A/n3563 , 
        \MAIN/ENGIN/STEP_A/n3561 , \MAIN/ENGIN/STEP_A/tmp2[2] , 
        \MAIN/ENGIN/STEP_A/n3571 , \MAIN/ENGIN/STEP_A/n3548 , 
        \MAIN/ENGIN/STEP_A/n3553 , \MAIN/ENGIN/STEP_A/n3554 , 
        \MAIN/ENGIN/STEP_A/n3584 , \MAIN/ENGIN/STEP_A/n3568 , 
        \MAIN/ENGIN/STEP_A/n3573 , \MAIN/ENGIN/STEP_A/n3574 , 
        \MAIN/ENGIN/STEP_A/n3566 , \MAIN/ENGIN/STEP_A/tmp2[1] , 
        \MAIN/ENGIN/STEP_A/n3583 , \MAIN/ENGIN/STEP_A/n3549 , 
        \MAIN/ENGIN/STEP_A/n3552 , \MAIN/ENGIN/STEP_A/n3590 , 
        \MAIN/ENGIN/STEP_A/n3567 , \MAIN/ENGIN/STEP_A/n3575 , 
        \MAIN/ENGIN/STEP_A/decode_stage272 , \MAIN/ENGIN/STEP_A/n3582 , 
        \MAIN/ENGIN/STEP_A/n3560 , \MAIN/ENGIN/STEP_A/n3585 , 
        \MAIN/ENGIN/STEP_A/n3547 , \MAIN/ENGIN/STEP_A/n3555 , 
        \MAIN/ENGIN/STEP_A/n3572 , \MAIN/ENGIN/STEP_A/d3_stage , 
        \MAIN/ENGIN/STEP_A/n3569 , \MAIN/ENGIN/STEP_B/cst[2] , 
        \MAIN/ENGIN/STEP_B/n3517 , \MAIN/ENGIN/STEP_B/n3530 , 
        \MAIN/ENGIN/STEP_B/n3505 , \MAIN/ENGIN/STEP_B/n3522 , 
        \MAIN/ENGIN/STEP_B/n3539 , \MAIN/ENGIN/STEP_B/n3519 , 
        \MAIN/ENGIN/STEP_B/cst[0] , \MAIN/ENGIN/STEP_B/n3502 , 
        \MAIN/ENGIN/STEP_B/n3525 , \MAIN/ENGIN/STEP_B/tmp2[0] , 
        \MAIN/ENGIN/STEP_B/n3510 , \MAIN/ENGIN/STEP_B/n3537 , 
        \MAIN/ENGIN/STEP_B/sw_stage , \MAIN/ENGIN/STEP_B/n3542 , 
        \MAIN/ENGIN/STEP_B/n3503 , \MAIN/ENGIN/STEP_B/n3524 , 
        \MAIN/ENGIN/STEP_B/nst[3] , \MAIN/ENGIN/STEP_B/cf_st2_rst , 
        \MAIN/ENGIN/STEP_B/n3511 , \MAIN/ENGIN/STEP_B/n3518 , 
        \MAIN/ENGIN/STEP_B/exec_stage278 , \MAIN/ENGIN/STEP_B/n3516 , 
        \MAIN/ENGIN/STEP_B/n3531 , \MAIN/ENGIN/STEP_B/n3536 , 
        \MAIN/ENGIN/STEP_B/cst[3] , \MAIN/ENGIN/STEP_B/cst[1] , 
        \MAIN/ENGIN/STEP_B/n3496 , \MAIN/ENGIN/STEP_B/n3504 , 
        \MAIN/ENGIN/STEP_B/dec_st2_rst , \MAIN/ENGIN/STEP_B/n3523 , 
        \MAIN/ENGIN/STEP_B/n3538 , \MAIN/ENGIN/STEP_B/n3506 , 
        \MAIN/ENGIN/STEP_B/n3514 , \MAIN/ENGIN/STEP_B/tmp2[2] , 
        \MAIN/ENGIN/STEP_B/n3528 , \MAIN/ENGIN/STEP_B/n3533 , 
        \MAIN/ENGIN/STEP_B/n3498 , \MAIN/ENGIN/STEP_B/n3501 , 
        \MAIN/ENGIN/STEP_B/n3521 , \MAIN/ENGIN/STEP_B/n3526 , 
        \MAIN/ENGIN/STEP_B/n3508 , \MAIN/ENGIN/STEP_B/n3513 , 
        \MAIN/ENGIN/STEP_B/n3534 , \MAIN/ENGIN/STEP_B/tmp2[1] , 
        \MAIN/ENGIN/STEP_B/n3541 , \MAIN/ENGIN/STEP_B/n3499 , 
        \MAIN/ENGIN/STEP_B/n3500 , \MAIN/ENGIN/STEP_B/n3527 , 
        \MAIN/ENGIN/STEP_B/n3540 , \MAIN/ENGIN/STEP_B/n3509 , 
        \MAIN/ENGIN/STEP_B/n3512 , \MAIN/ENGIN/STEP_B/decode_stage272 , 
        \MAIN/ENGIN/STEP_B/n3535 , \MAIN/ENGIN/STEP_B/n3515 , 
        \MAIN/ENGIN/STEP_B/n3529 , \MAIN/ENGIN/STEP_B/n3532 , 
        \MAIN/ENGIN/STEP_B/n3497 , \MAIN/ENGIN/STEP_B/d3_stage , 
        \MAIN/ENGIN/STEP_B/n3507 , \MAIN/ENGIN/STEP_B/n3520 , 
        \MAIN/ENGIN/STEP_C/cst[2] , \MAIN/ENGIN/STEP_C/n3462 , 
        \MAIN/ENGIN/STEP_C/n3479 , \MAIN/ENGIN/STEP_C/n3487 , 
        \MAIN/ENGIN/STEP_C/n3457 , \MAIN/ENGIN/STEP_C/n3470 , 
        \MAIN/ENGIN/STEP_C/n3489 , \MAIN/ENGIN/STEP_C/cst[0] , 
        \MAIN/ENGIN/STEP_C/n3450 , \MAIN/ENGIN/STEP_C/n3492 , 
        \MAIN/ENGIN/STEP_C/n3465 , \MAIN/ENGIN/STEP_C/n3477 , 
        \MAIN/ENGIN/STEP_C/tmp2[0] , \MAIN/ENGIN/STEP_C/n3459 , 
        \MAIN/ENGIN/STEP_C/n3480 , \MAIN/ENGIN/STEP_C/sw_stage , 
        \MAIN/ENGIN/STEP_C/n3451 , \MAIN/ENGIN/STEP_C/n3476 , 
        \MAIN/ENGIN/STEP_C/n3493 , \MAIN/ENGIN/STEP_C/n3458 , 
        \MAIN/ENGIN/STEP_C/nst[3] , \MAIN/ENGIN/STEP_C/exec_stage278 , 
        \MAIN/ENGIN/STEP_C/n3488 , \MAIN/ENGIN/STEP_C/cf_st2_rst , 
        \MAIN/ENGIN/STEP_C/n3481 , \MAIN/ENGIN/STEP_C/n3463 , 
        \MAIN/ENGIN/STEP_C/n3464 , \MAIN/ENGIN/STEP_C/n3486 , 
        \MAIN/ENGIN/STEP_C/cst[3] , \MAIN/ENGIN/STEP_C/cst[1] , 
        \MAIN/ENGIN/STEP_C/n3448 , \MAIN/ENGIN/STEP_C/n3454 , 
        \MAIN/ENGIN/STEP_C/n3456 , \MAIN/ENGIN/STEP_C/dec_st2_rst , 
        \MAIN/ENGIN/STEP_C/n3471 , \MAIN/ENGIN/STEP_C/tmp2[2] , 
        \MAIN/ENGIN/STEP_C/n3478 , \MAIN/ENGIN/STEP_C/n3494 , 
        \MAIN/ENGIN/STEP_C/n3461 , \MAIN/ENGIN/STEP_C/n3484 , 
        \MAIN/ENGIN/STEP_C/n3468 , \MAIN/ENGIN/STEP_C/n3473 , 
        \MAIN/ENGIN/STEP_C/n3452 , \MAIN/ENGIN/STEP_C/n3453 , 
        \MAIN/ENGIN/STEP_C/n3474 , \MAIN/ENGIN/STEP_C/n3491 , 
        \MAIN/ENGIN/STEP_C/n3466 , \MAIN/ENGIN/STEP_C/n3483 , 
        \MAIN/ENGIN/STEP_C/tmp2[1] , \MAIN/ENGIN/STEP_C/n3475 , 
        \MAIN/ENGIN/STEP_C/n3449 , \MAIN/ENGIN/STEP_C/n3490 , 
        \MAIN/ENGIN/STEP_C/n3460 , \MAIN/ENGIN/STEP_C/decode_stage272 , 
        \MAIN/ENGIN/STEP_C/n3467 , \MAIN/ENGIN/STEP_C/n3482 , 
        \MAIN/ENGIN/STEP_C/n3485 , \MAIN/ENGIN/STEP_C/n3455 , 
        \MAIN/ENGIN/STEP_C/n3469 , \MAIN/ENGIN/STEP_C/d3_stage , 
        \MAIN/ENGIN/STEP_C/n3472 , \MAIN/ENGIN/STEP_D/cst[2] , 
        \MAIN/ENGIN/STEP_D/n3417 , \MAIN/ENGIN/STEP_D/n3430 , 
        \MAIN/ENGIN/STEP_D/n3445 , \MAIN/ENGIN/STEP_D/n3405 , 
        \MAIN/ENGIN/STEP_D/n3439 , \MAIN/ENGIN/STEP_D/n3422 , 
        \MAIN/ENGIN/STEP_D/cst[0] , \MAIN/ENGIN/STEP_D/n3402 , 
        \MAIN/ENGIN/STEP_D/n3425 , \MAIN/ENGIN/STEP_D/n3419 , 
        \MAIN/ENGIN/STEP_D/n3442 , \MAIN/ENGIN/STEP_D/tmp2[0] , 
        \MAIN/ENGIN/STEP_D/n3410 , \MAIN/ENGIN/STEP_D/n3437 , 
        \MAIN/ENGIN/STEP_D/sw_stage , \MAIN/ENGIN/STEP_D/n3403 , 
        \MAIN/ENGIN/STEP_D/n3418 , \MAIN/ENGIN/STEP_D/nst[3] , 
        \MAIN/ENGIN/STEP_D/exec_stage278 , \MAIN/ENGIN/STEP_D/n3424 , 
        \MAIN/ENGIN/STEP_D/n3411 , \MAIN/ENGIN/STEP_D/n3436 , 
        \MAIN/ENGIN/STEP_D/cf_st2_rst , \MAIN/ENGIN/STEP_D/n3416 , 
        \MAIN/ENGIN/STEP_D/n3443 , \MAIN/ENGIN/STEP_D/n3444 , 
        \MAIN/ENGIN/STEP_D/cst[3] , \MAIN/ENGIN/STEP_D/cst[1] , 
        \MAIN/ENGIN/STEP_D/n3401 , \MAIN/ENGIN/STEP_D/n3404 , 
        \MAIN/ENGIN/STEP_D/dec_st2_rst , \MAIN/ENGIN/STEP_D/n3431 , 
        \MAIN/ENGIN/STEP_D/n3406 , \MAIN/ENGIN/STEP_D/n3414 , 
        \MAIN/ENGIN/STEP_D/n3423 , \MAIN/ENGIN/STEP_D/tmp2[2] , 
        \MAIN/ENGIN/STEP_D/n3438 , \MAIN/ENGIN/STEP_D/n3433 , 
        \MAIN/ENGIN/STEP_D/n3428 , \MAIN/ENGIN/STEP_D/n3446 , 
        \MAIN/ENGIN/STEP_D/n3421 , \MAIN/ENGIN/STEP_D/n3408 , 
        \MAIN/ENGIN/STEP_D/n3426 , \MAIN/ENGIN/STEP_D/n3441 , 
        \MAIN/ENGIN/STEP_D/tmp2[1] , \MAIN/ENGIN/STEP_D/n3413 , 
        \MAIN/ENGIN/STEP_D/n3434 , \MAIN/ENGIN/STEP_D/n3400 , 
        \MAIN/ENGIN/STEP_D/n3409 , \MAIN/ENGIN/STEP_D/n3412 , 
        \MAIN/ENGIN/STEP_D/n3427 , \MAIN/ENGIN/STEP_D/n3435 , 
        \MAIN/ENGIN/STEP_D/decode_stage272 , \MAIN/ENGIN/STEP_D/n3440 , 
        \MAIN/ENGIN/STEP_D/n3415 , \MAIN/ENGIN/STEP_D/n3429 , 
        \MAIN/ENGIN/STEP_D/n3432 , \MAIN/ENGIN/STEP_D/n3407 , 
        \MAIN/ENGIN/STEP_D/n3420 , \MAIN/ENGIN/STEP_D/d3_stage , 
        \CONS/phinc20_1/inc4_1/n325 , \CONS/phinc20_1/inc4_1/n326 , 
        \CONS/phinc20_1/inc4_1/n327 , \CONS/phinc20_1/inc4_2/n322 , 
        \CONS/phinc20_1/inc4_2/n324 , \CONS/phinc20_1/inc4_2/n323 , 
        \CONS/phinc20_1/inc4_3/n319 , \CONS/phinc20_1/inc4_3/n321 , 
        \CONS/phinc20_1/inc4_3/n320 , \CONS/phinc20_1/inc4_4/n317 , 
        \CONS/phinc20_1/inc4_4/n316 , \CONS/phinc20_1/inc4_4/n318 , 
        \CONS/phinc20_1/inc4_5/gp_out , \CONS/phinc20_1/inc4_5/n311 , 
        \CONS/phinc20_1/inc4_5/n312 , \CONS/phinc20_1/inc4_5/n313 , 
        \CONS/phinc20_1/inc4_5/n314 , \CONS/phinc20_1/inc4_5/n315 , 
        \CODEIF/inc19_1/inc4_1/n3760 , \CODEIF/inc19_1/inc4_1/n3761 , 
        \CODEIF/inc19_1/inc4_1/n3762 , \CODEIF/inc19_1/inc4_2/n3758 , 
        \CODEIF/inc19_1/inc4_2/n3757 , \CODEIF/inc19_1/inc4_2/n3759 , 
        \CODEIF/inc19_1/inc4_3/n3755 , \CODEIF/inc19_1/inc4_3/n3656 , 
        \CODEIF/inc19_1/inc4_3/n3756 , \CODEIF/inc19_1/inc4_4/n3652 , 
        \CODEIF/inc19_1/inc4_4/n3654 , \CODEIF/inc19_1/inc4_4/n3650 , 
        \CODEIF/inc19_1/inc4_5/gp_out , \CODEIF/inc19_1/inc4_5/n3640 , 
        \CODEIF/inc19_1/inc4_5/n3646 , \CODEIF/inc19_1/inc4_5/n3648 , 
        \CODEIF/inc19_1/inc4_5/n3644 , \CODEIF/inc19_1/inc4_5/n3642 , 
        \UPIF/RCTL/regfile_1/n1020 , \UPIF/RCTL/regfile_1/n1021 , 
        \UPIF/RCTL/regfile_1/n1016 , \UPIF/RCTL/regfile_1/n1018 , 
        \UPIF/RCTL/regfile_1/n1019 , \UPIF/RCTL/regfile_1/n1017 , 
        \UPIF/RCTL/regfile_1/n1022 , 
        \REGF/pbmemff31/SACNST/*cell*5426/U1/CONTROL2 , 
        \REGF/pbmemff31/SACNST/n5645 , \REGF/pbmemff31/SACNST/n5646 , 
        \ALUSHT/ALU/dec32/gg_out[4] , \ALUSHT/ALU/dec32/gg_out[0] , 
        \ALUSHT/ALU/dec32/gg_out[2] , \ALUSHT/ALU/dec32/gg_out[6] , 
        \ALUSHT/ALU/dec32/n1801 , \ALUSHT/ALU/dec32/gcarry[1] , 
        \ALUSHT/ALU/dec32/gcarry[5] , \ALUSHT/ALU/dec32/gcarry[3] , 
        \ALUSHT/ALU/dec32/gcarry[2] , \ALUSHT/ALU/dec32/gcarry[6] , 
        \ALUSHT/ALU/dec32/gcarry[4] , \ALUSHT/ALU/dec32/gg_out[1] , 
        \ALUSHT/ALU/dec32/gg_out[3] , \ALUSHT/ALU/dec32/gg_out[5] , 
        \ALUSHT/ALU/add32/gg_out[0] , \ALUSHT/ALU/add32/gg_out[4] , 
        \ALUSHT/ALU/add32/c_last , \ALUSHT/ALU/add32/n1389 , 
        \ALUSHT/ALU/add32/gg_out[2] , \ALUSHT/ALU/add32/n1394 , 
        \ALUSHT/ALU/add32/gp_out[3] , \ALUSHT/ALU/add32/cin_stg[3] , 
        \ALUSHT/ALU/add32/cin_stg[1] , \ALUSHT/ALU/add32/gp_out[5] , 
        \ALUSHT/ALU/add32/gp_out[1] , \ALUSHT/ALU/add32/cin_stg[4] , 
        \ALUSHT/ALU/add32/gp_out[0] , \ALUSHT/ALU/add32/cin_stg[0] , 
        \ALUSHT/ALU/add32/gp_out[4] , \ALUSHT/ALU/add32/cin_stg[2] , 
        \ALUSHT/ALU/add32/gp_out[2] , \ALUSHT/ALU/add32/n1635 , 
        \ALUSHT/ALU/add32/gg_out[1] , \ALUSHT/ALU/add32/gg_out[3] , 
        \ALUSHT/ALU/add32/gg_out[5] , \ALUSHT/ALU/add32/n1390 , 
        \ALUSHT/ALU/cmp32/ggflg[7] , \ALUSHT/ALU/cmp32/geqflg[0] , 
        \ALUSHT/ALU/cmp32/ggflg[6] , \ALUSHT/ALU/cmp32/geqflg[4] , 
        \ALUSHT/ALU/cmp32/ggflg[0] , \ALUSHT/ALU/cmp32/ggflg[2] , 
        \ALUSHT/ALU/cmp32/n1219 , \ALUSHT/ALU/cmp32/geqflg[7] , 
        \ALUSHT/ALU/cmp32/geqflg[6] , \ALUSHT/ALU/cmp32/n1217 , 
        \ALUSHT/ALU/cmp32/ggflg[4] , \ALUSHT/ALU/cmp32/geqflg[2] , 
        \ALUSHT/ALU/cmp32/n1216 , \ALUSHT/ALU/cmp32/n1211 , 
        \ALUSHT/ALU/cmp32/n1218 , \ALUSHT/ALU/cmp32/n1213 , 
        \ALUSHT/ALU/cmp32/n1214 , \ALUSHT/ALU/cmp32/n1220 , 
        \ALUSHT/ALU/cmp32/ggflg[5] , \ALUSHT/ALU/cmp32/geqflg[3] , 
        \ALUSHT/ALU/cmp32/ggflg[1] , \ALUSHT/ALU/cmp32/n1212 , 
        \ALUSHT/ALU/cmp32/n1215 , \ALUSHT/ALU/cmp32/geqflg[5] , 
        \ALUSHT/ALU/cmp32/geqflg[1] , \ALUSHT/ALU/cmp32/ggflg[3] , 
        \ALUSHT/ALU/inc32/gg_out[4] , \ALUSHT/ALU/inc32/gg_out[2] , 
        \ALUSHT/ALU/inc32/gg_out[6] , \ALUSHT/ALU/inc32/gp_out[3] , 
        \ALUSHT/ALU/inc32/gp_out[5] , \ALUSHT/ALU/inc32/gp_out[1] , 
        \ALUSHT/ALU/inc32/gp_out[0] , \ALUSHT/ALU/inc32/gp_out[6] , 
        \ALUSHT/ALU/inc32/gp_out[4] , \ALUSHT/ALU/inc32/gp_out[2] , 
        \ALUSHT/ALU/inc32/gg_out[1] , \ALUSHT/ALU/inc32/gg_out[3] , 
        \ALUSHT/ALU/inc32/gg_out[5] , \MAIN/STM/SEQMG/n3346 , 
        \MAIN/STM/SEQMG/n3354 , \MAIN/STM/SEQMG/eqst[0] , 
        \MAIN/STM/SEQMG/n3361 , \MAIN/STM/SEQMG/n3348 , \MAIN/STM/SEQMG/n3353 , 
        \MAIN/STM/SEQMG/n3345 , \MAIN/STM/SEQMG/n3347 , \MAIN/STM/SEQMG/n3349 , 
        \MAIN/STM/SEQMG/n3352 , \MAIN/STM/SEQMG/n3355 , \MAIN/STM/SEQMG/n3357 , 
        \MAIN/STM/SEQMG/n3360 , \MAIN/STM/SEQMG/n3362 , \MAIN/STM/SEQMG/n3350 , 
        \MAIN/STM/SEQMG/n3359 , \MAIN/STM/SEQMG/n3351 , \MAIN/STM/SEQMG/n3358 , 
        \MAIN/STM/SEQMG/temp[1] , \MAIN/STM/SEQMG/n3356 , 
        \MAIN/STM/SEQMG/eqst[1] , \MAIN/STM/NS/n3341 , \MAIN/STM/NS/n3338 , 
        \MAIN/STM/NS/est[1] , \MAIN/STM/NS/n3339 , \MAIN/STM/NS/n3340 , 
        \MAIN/STM/NS/nst[0] , \MAIN/STM/NS/nst[1] , \MAIN/STM/NS/n3342 , 
        \MAIN/STM/NS/n3343 , \MAIN/STM/NS/n3344 , \MAIN/STM/WS/nwst[1] , 
        \MAIN/STM/WS/ewst[0] , \MAIN/STM/WS/n3333 , \MAIN/STM/WS/n3334 , 
        \MAIN/STM/WS/n3335 , \MAIN/STM/WS/n3336 , \MAIN/STM/WS/n3337 , 
        \MAIN/STM/WS/ewst[1] , \MAIN/STM/RS/n3328 , \MAIN/STM/RS/nrst[0] , 
        \MAIN/STM/RS/n3326 , \MAIN/STM/RS/n3327 , \MAIN/STM/RS/n3324 , 
        \MAIN/STM/RS/n3325 , \MAIN/STM/RS/n3329 , \MAIN/STM/RS/erst[1] , 
        \MAIN/STM/RS/n3332 , \MAIN/STM/RS/n3330 , \MAIN/STM/RS/erst[0] , 
        \MAIN/STM/RS/n3331 , \SAEXE/RFIO/phcont4_1/ph4dec_1/n14 , 
        \SADR/MAINSADR/addidxof/add0/c_last , 
        \SADR/MAINSADR/addidxof/add0/n8607 , 
        \SADR/MAINSADR/addidxof/add0/n8620 , 
        \SADR/MAINSADR/addidxof/add0/n8629 , 
        \SADR/MAINSADR/addidxof/add0/n8612 , 
        \SADR/MAINSADR/addidxof/add0/n8615 , 
        \SADR/MAINSADR/addidxof/add0/n8600 , 
        \SADR/MAINSADR/addidxof/add0/n8609 , 
        \SADR/MAINSADR/addidxof/add0/n8601 , 
        \SADR/MAINSADR/addidxof/add0/n8608 , 
        \SADR/MAINSADR/addidxof/add0/n8627 , 
        \SADR/MAINSADR/addidxof/add0/n8613 , 
        \SADR/MAINSADR/addidxof/add0/n8602 , 
        \SADR/MAINSADR/addidxof/add0/gp_out , 
        \SADR/MAINSADR/addidxof/add0/n8606 , 
        \SADR/MAINSADR/addidxof/add0/n8621 , 
        \SADR/MAINSADR/addidxof/add0/n8626 , 
        \SADR/MAINSADR/addidxof/add0/n8614 , 
        \SADR/MAINSADR/addidxof/add0/n8603 , 
        \SADR/MAINSADR/addidxof/add0/n8604 , 
        \SADR/MAINSADR/addidxof/add0/n8628 , 
        \SADR/MAINSADR/addidxof/add0/n8611 , 
        \SADR/MAINSADR/addidxof/add0/n8616 , 
        \SADR/MAINSADR/addidxof/add0/n8623 , 
        \SADR/MAINSADR/addidxof/add0/n8631 , 
        \SADR/MAINSADR/addidxof/add0/n8618 , 
        \SADR/MAINSADR/addidxof/add0/n8624 , 
        \SADR/MAINSADR/addidxof/add0/n8610 , 
        \SADR/MAINSADR/addidxof/add0/n8625 , 
        \SADR/MAINSADR/addidxof/add0/n8605 , 
        \SADR/MAINSADR/addidxof/add0/n8619 , 
        \SADR/MAINSADR/addidxof/add0/n8617 , 
        \SADR/MAINSADR/addidxof/add0/n8622 , 
        \SADR/MAINSADR/addidxof/add0/n8630 , 
        \SADR/MAINSADR/addidxof/add1/c_last , 
        \SADR/MAINSADR/addidxof/add1/n8577 , 
        \SADR/MAINSADR/addidxof/add1/n8580 , 
        \SADR/MAINSADR/addidxof/add1/n8592 , 
        \SADR/MAINSADR/addidxof/add1/n8589 , 
        \SADR/MAINSADR/addidxof/add1/n8568 , 
        \SADR/MAINSADR/addidxof/add1/n8570 , 
        \SADR/MAINSADR/addidxof/add1/n8571 , 
        \SADR/MAINSADR/addidxof/add1/n8579 , 
        \SADR/MAINSADR/addidxof/add1/n8587 , 
        \SADR/MAINSADR/addidxof/add1/n8595 , 
        \SADR/MAINSADR/addidxof/add1/n8594 , 
        \SADR/MAINSADR/addidxof/add1/n8578 , 
        \SADR/MAINSADR/addidxof/add1/n8581 , 
        \SADR/MAINSADR/addidxof/add1/n8586 , 
        \SADR/MAINSADR/addidxof/add1/n8588 , 
        \SADR/MAINSADR/addidxof/add1/n8574 , 
        \SADR/MAINSADR/addidxof/add1/n8576 , 
        \SADR/MAINSADR/addidxof/add1/n8593 , 
        \SADR/MAINSADR/addidxof/add1/n8583 , 
        \SADR/MAINSADR/addidxof/add1/n8598 , 
        \SADR/MAINSADR/addidxof/add1/n8591 , 
        \SADR/MAINSADR/addidxof/add1/n8569 , 
        \SADR/MAINSADR/addidxof/add1/n8572 , 
        \SADR/MAINSADR/addidxof/add1/n8573 , 
        \SADR/MAINSADR/addidxof/add1/n8584 , 
        \SADR/MAINSADR/addidxof/add1/n8596 , 
        \SADR/MAINSADR/addidxof/add1/n8597 , 
        \SADR/MAINSADR/addidxof/add1/n8575 , 
        \SADR/MAINSADR/addidxof/add1/n8582 , 
        \SADR/MAINSADR/addidxof/add1/n8585 , 
        \SADR/MAINSADR/addidxof/add1/n8599 , 
        \SADR/MAINSADR/addidxof/add1/n8590 , 
        \SADR/MAINSADR/addidxof/add2/c_last , 
        \SADR/MAINSADR/addidxof/add2/n8537 , 
        \SADR/MAINSADR/addidxof/add2/n8542 , 
        \SADR/MAINSADR/addidxof/add2/n8559 , 
        \SADR/MAINSADR/addidxof/add2/n8565 , 
        \SADR/MAINSADR/addidxof/add2/n8550 , 
        \SADR/MAINSADR/addidxof/add2/n8536 , 
        \SADR/MAINSADR/addidxof/add2/n8538 , 
        \SADR/MAINSADR/addidxof/add2/n8539 , 
        \SADR/MAINSADR/addidxof/add2/n8557 , 
        \SADR/MAINSADR/addidxof/add2/n8545 , 
        \SADR/MAINSADR/addidxof/add2/n8562 , 
        \SADR/MAINSADR/addidxof/add2/n8543 , 
        \SADR/MAINSADR/addidxof/add2/n8544 , 
        \SADR/MAINSADR/addidxof/add2/n8556 , 
        \SADR/MAINSADR/addidxof/add2/n8563 , 
        \SADR/MAINSADR/addidxof/add2/n8564 , 
        \SADR/MAINSADR/addidxof/add2/n8558 , 
        \SADR/MAINSADR/addidxof/add2/n8540 , 
        \SADR/MAINSADR/addidxof/add2/n8541 , 
        \SADR/MAINSADR/addidxof/add2/n8551 , 
        \SADR/MAINSADR/addidxof/add2/n8546 , 
        \SADR/MAINSADR/addidxof/add2/n8548 , 
        \SADR/MAINSADR/addidxof/add2/n8553 , 
        \SADR/MAINSADR/addidxof/add2/n8566 , 
        \SADR/MAINSADR/addidxof/add2/n8554 , 
        \SADR/MAINSADR/addidxof/add2/n8561 , 
        \SADR/MAINSADR/addidxof/add2/n8547 , 
        \SADR/MAINSADR/addidxof/add2/n8555 , 
        \SADR/MAINSADR/addidxof/add2/n8560 , 
        \SADR/MAINSADR/addidxof/add2/n8549 , 
        \SADR/MAINSADR/addidxof/add2/n8567 , 
        \SADR/MAINSADR/addidxof/add2/n8552 , 
        \SADR/MAINSADR/addidxof/add3/n8510 , 
        \SADR/MAINSADR/addidxof/add3/n8519 , 
        \SADR/MAINSADR/addidxof/add3/n8505 , 
        \SADR/MAINSADR/addidxof/add3/n8522 , 
        \SADR/MAINSADR/addidxof/add3/n8525 , 
        \SADR/MAINSADR/addidxof/add3/n8504 , 
        \SADR/MAINSADR/addidxof/add3/n8517 , 
        \SADR/MAINSADR/addidxof/add3/n8530 , 
        \SADR/MAINSADR/addidxof/add3/n8523 , 
        \SADR/MAINSADR/addidxof/add3/n8506 , 
        \SADR/MAINSADR/addidxof/add3/n8511 , 
        \SADR/MAINSADR/addidxof/add3/n8516 , 
        \SADR/MAINSADR/addidxof/add3/n8531 , 
        \SADR/MAINSADR/addidxof/add3/n8524 , 
        \SADR/MAINSADR/addidxof/add3/n8508 , 
        \SADR/MAINSADR/addidxof/add3/n8513 , 
        \SADR/MAINSADR/addidxof/add3/n8518 , 
        \SADR/MAINSADR/addidxof/add3/n8534 , 
        \SADR/MAINSADR/addidxof/add3/n8526 , 
        \SADR/MAINSADR/addidxof/add3/n8507 , 
        \SADR/MAINSADR/addidxof/add3/n8514 , 
        \SADR/MAINSADR/addidxof/add3/n8521 , 
        \SADR/MAINSADR/addidxof/add3/n8528 , 
        \SADR/MAINSADR/addidxof/add3/n8533 , 
        \SADR/MAINSADR/addidxof/add3/n8509 , 
        \SADR/MAINSADR/addidxof/add3/n8515 , 
        \SADR/MAINSADR/addidxof/add3/n8520 , 
        \SADR/MAINSADR/addidxof/add3/n8532 , 
        \SADR/MAINSADR/addidxof/add3/n8529 , 
        \SADR/MAINSADR/addidxof/add3/n8512 , 
        \SADR/MAINSADR/addidxof/add3/n8535 , 
        \SADR/MAINSADR/addidxof/add3/n8527 , 
        \SADR/MAINSADR/addsegoff/add0/gp_out , 
        \SADR/MAINSADR/addsegoff/add0/n8465 , 
        \SADR/MAINSADR/addsegoff/add0/n8480 , 
        \SADR/MAINSADR/addsegoff/add0/n8470 , 
        \SADR/MAINSADR/addsegoff/add0/n8477 , 
        \SADR/MAINSADR/addsegoff/add0/n8489 , 
        \SADR/MAINSADR/addsegoff/add0/n8492 , 
        \SADR/MAINSADR/addsegoff/add0/n8495 , 
        \SADR/MAINSADR/addsegoff/add0/n8462 , 
        \SADR/MAINSADR/addsegoff/add0/n8479 , 
        \SADR/MAINSADR/addsegoff/add0/n8463 , 
        \SADR/MAINSADR/addsegoff/add0/n8471 , 
        \SADR/MAINSADR/addsegoff/add0/n8487 , 
        \SADR/MAINSADR/addsegoff/add0/n8486 , 
        \SADR/MAINSADR/addsegoff/add0/n8494 , 
        \SADR/MAINSADR/addsegoff/add0/n8464 , 
        \SADR/MAINSADR/addsegoff/add0/n8478 , 
        \SADR/MAINSADR/addsegoff/add0/n8481 , 
        \SADR/MAINSADR/addsegoff/add0/n8493 , 
        \SADR/MAINSADR/addsegoff/add0/n8461 , 
        \SADR/MAINSADR/addsegoff/add0/n8476 , 
        \SADR/MAINSADR/addsegoff/add0/n8466 , 
        \SADR/MAINSADR/addsegoff/add0/n8483 , 
        \SADR/MAINSADR/addsegoff/add0/n8488 , 
        \SADR/MAINSADR/addsegoff/add0/n8468 , 
        \SADR/MAINSADR/addsegoff/add0/n8473 , 
        \SADR/MAINSADR/addsegoff/add0/n8474 , 
        \SADR/MAINSADR/addsegoff/add0/n8491 , 
        \SADR/MAINSADR/addsegoff/add0/n8496 , 
        \SADR/MAINSADR/addsegoff/add0/n8467 , 
        \SADR/MAINSADR/addsegoff/add0/n8469 , 
        \SADR/MAINSADR/addsegoff/add0/n8484 , 
        \SADR/MAINSADR/addsegoff/add0/n8472 , 
        \SADR/MAINSADR/addsegoff/add0/n8485 , 
        \SADR/MAINSADR/addsegoff/add0/n8475 , 
        \SADR/MAINSADR/addsegoff/add0/n8482 , 
        \SADR/MAINSADR/addsegoff/add0/n8490 , 
        \SADR/MAINSADR/addsegoff/add1/n8425 , 
        \SADR/MAINSADR/addsegoff/add1/n8437 , 
        \SADR/MAINSADR/addsegoff/add1/n8442 , 
        \SADR/MAINSADR/addsegoff/add1/n8459 , 
        \SADR/MAINSADR/addsegoff/add1/n8439 , 
        \SADR/MAINSADR/addsegoff/add1/n8450 , 
        \SADR/MAINSADR/addsegoff/add1/n8457 , 
        \SADR/MAINSADR/addsegoff/add1/n8430 , 
        \SADR/MAINSADR/addsegoff/add1/n8431 , 
        \SADR/MAINSADR/addsegoff/add1/n8438 , 
        \SADR/MAINSADR/addsegoff/add1/n8445 , 
        \SADR/MAINSADR/addsegoff/add1/n8456 , 
        \SADR/MAINSADR/addsegoff/add1/n8444 , 
        \SADR/MAINSADR/addsegoff/add1/n8436 , 
        \SADR/MAINSADR/addsegoff/add1/n8443 , 
        \SADR/MAINSADR/addsegoff/add1/n8458 , 
        \SADR/MAINSADR/addsegoff/add1/n8426 , 
        \SADR/MAINSADR/addsegoff/add1/n8451 , 
        \SADR/MAINSADR/addsegoff/add1/n8434 , 
        \SADR/MAINSADR/addsegoff/add1/n8441 , 
        \SADR/MAINSADR/addsegoff/add1/n8427 , 
        \SADR/MAINSADR/addsegoff/add1/n8428 , 
        \SADR/MAINSADR/addsegoff/add1/n8433 , 
        \SADR/MAINSADR/addsegoff/add1/n8448 , 
        \SADR/MAINSADR/addsegoff/add1/n8453 , 
        \SADR/MAINSADR/addsegoff/add1/n8454 , 
        \SADR/MAINSADR/addsegoff/add1/n8446 , 
        \SADR/MAINSADR/addsegoff/add1/n8429 , 
        \SADR/MAINSADR/addsegoff/add1/n8455 , 
        \SADR/MAINSADR/addsegoff/add1/n8432 , 
        \SADR/MAINSADR/addsegoff/add1/n8447 , 
        \SADR/MAINSADR/addsegoff/add1/n8460 , 
        \SADR/MAINSADR/addsegoff/add1/n8435 , 
        \SADR/MAINSADR/addsegoff/add1/n8440 , 
        \SADR/MAINSADR/addsegoff/add1/n8449 , 
        \SADR/MAINSADR/addsegoff/add1/n8452 , 
        \SADR/MAINSADR/adrinc1/inc4_1/n8422 , 
        \SADR/MAINSADR/adrinc1/inc4_1/n8423 , 
        \SADR/MAINSADR/adrinc1/inc4_1/n8424 , 
        \SADR/MAINSADR/adrinc1/inc4_6/gp_out , 
        \SADR/MAINSADR/adrinc1/inc4_6/n8419 , 
        \SADR/MAINSADR/adrinc1/inc4_6/n8420 , 
        \SADR/MAINSADR/adrinc1/inc4_6/n8421 , 
        \SADR/MAINSADR/adrinc1/inc4_2/n8416 , 
        \SADR/MAINSADR/adrinc1/inc4_2/n8417 , 
        \SADR/MAINSADR/adrinc1/inc4_2/n8418 , 
        \SADR/MAINSADR/adrinc1/inc4_3/n8413 , 
        \SADR/MAINSADR/adrinc1/inc4_3/n8414 , 
        \SADR/MAINSADR/adrinc1/inc4_3/n8415 , 
        \SADR/MAINSADR/adrinc1/inc4_4/n8410 , 
        \SADR/MAINSADR/adrinc1/inc4_4/n8411 , 
        \SADR/MAINSADR/adrinc1/inc4_4/n8412 , 
        \SADR/MAINSADR/adrinc1/inc4_5/n8407 , 
        \SADR/MAINSADR/adrinc1/inc4_5/n8408 , 
        \SADR/MAINSADR/adrinc1/inc4_5/n8409 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8391 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8402 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8398 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8396 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8390 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8397 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8392 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8399 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8403 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8395 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8401 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8393 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8394 , 
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8400 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8383 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8384 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8377 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8382 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8385 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8389 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8378 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8379 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8380 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8386 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8387 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8376 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8381 , 
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8388 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8366 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8374 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8362 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8365 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8367 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8368 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8373 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8369 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8372 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8375 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8363 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8370 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8371 , 
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8364 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8348 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8353 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8361 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8349 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8352 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8354 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8355 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8360 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8350 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8357 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8359 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8351 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8356 , 
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8358 , 
        \SADR/MAINSADR/adrdec1/dec4_1/n8346 , 
        \SADR/MAINSADR/adrdec1/dec4_1/n8342 , 
        \SADR/MAINSADR/adrdec1/dec4_1/n8345 , 
        \SADR/MAINSADR/adrdec1/dec4_1/n8344 , 
        \SADR/MAINSADR/adrdec1/dec4_1/n8343 , 
        \SADR/MAINSADR/adrdec1/dec4_2/n8341 , 
        \SADR/MAINSADR/adrdec1/dec4_2/n8340 , 
        \SADR/MAINSADR/adrdec1/dec4_2/n8337 , 
        \SADR/MAINSADR/adrdec1/dec4_2/n8339 , 
        \SADR/MAINSADR/adrdec1/dec4_2/n8338 , 
        \SADR/MAINSADR/adrdec1/dec4_3/n8333 , 
        \SADR/MAINSADR/adrdec1/dec4_3/n8334 , 
        \SADR/MAINSADR/adrdec1/dec4_3/n8332 , 
        \SADR/MAINSADR/adrdec1/dec4_3/n8335 , 
        \SADR/MAINSADR/adrdec1/dec4_3/n8336 , 
        \SADR/MAINSADR/adrdec1/dec4_4/n8328 , 
        \SADR/MAINSADR/adrdec1/dec4_4/n8329 , 
        \SADR/MAINSADR/adrdec1/dec4_4/n8327 , 
        \SADR/MAINSADR/adrdec1/dec4_4/n8330 , 
        \SADR/MAINSADR/adrdec1/dec4_4/n8331 , 
        \SADR/MAINSADR/adrdec1/dec4_6/n8326 , 
        \SADR/MAINSADR/adrdec1/dec4_6/gg_out , 
        \SADR/MAINSADR/adrdec1/dec4_6/n8325 , 
        \SADR/MAINSADR/adrdec1/dec4_6/n8322 , 
        \SADR/MAINSADR/adrdec1/dec4_6/n8323 , 
        \SADR/MAINSADR/adrdec1/dec4_6/n8324 , 
        \SADR/MAINSADR/adrdec1/dec4_5/n8321 , 
        \SADR/MAINSADR/adrdec1/dec4_5/n8320 , 
        \SADR/MAINSADR/adrdec1/dec4_5/n8317 , 
        \SADR/MAINSADR/adrdec1/dec4_5/n8319 , 
        \SADR/MAINSADR/adrdec1/dec4_5/n8318 , 
        \SADR/MAINSADR/adrinc2/inc4_1/n8314 , 
        \SADR/MAINSADR/adrinc2/inc4_1/n8315 , 
        \SADR/MAINSADR/adrinc2/inc4_1/n8316 , 
        \SADR/MAINSADR/adrinc2/inc4_2/n8313 , 
        \SADR/MAINSADR/adrinc2/inc4_2/n8312 , 
        \SADR/MAINSADR/adrinc2/inc4_2/n8311 , 
        \SADR/MAINSADR/adrinc2/inc4_3/n8308 , 
        \SADR/MAINSADR/adrinc2/inc4_3/n8309 , 
        \SADR/MAINSADR/adrinc2/inc4_3/n8310 , 
        \SADR/MAINSADR/adrinc2/inc4_4/n8306 , 
        \SADR/MAINSADR/adrinc2/inc4_4/n8307 , 
        \SADR/MAINSADR/adrinc2/inc4_4/n8305 , 
        \SADR/MAINSADR/adrinc2/inc4_5/n8302 , 
        \SADR/MAINSADR/adrinc2/inc4_5/n8304 , 
        \SADR/MAINSADR/adrinc2/inc4_5/n8303 , 
        \SADR/MAINSADR/adrinc2/inc3_6/gp_out , 
        \SADR/MAINSADR/adrinc2/inc3_6/n8301 , 
        \SADR/MAINSADR/adrinc2/inc3_6/n8300 , 
        \SADR/MAINSADR/adrdec2/dec4_1/n8298 , 
        \SADR/MAINSADR/adrdec2/dec4_1/n8296 , 
        \SADR/MAINSADR/adrdec2/dec4_1/n8297 , 
        \SADR/MAINSADR/adrdec2/dec4_1/n8294 , 
        \SADR/MAINSADR/adrdec2/dec4_1/n8295 , 
        \SADR/MAINSADR/adrdec2/dec4_2/n8291 , 
        \SADR/MAINSADR/adrdec2/dec4_2/n8290 , 
        \SADR/MAINSADR/adrdec2/dec4_2/n8292 , 
        \SADR/MAINSADR/adrdec2/dec4_2/n8289 , 
        \SADR/MAINSADR/adrdec2/dec4_2/n8293 , 
        \SADR/MAINSADR/adrdec2/dec4_3/n8284 , 
        \SADR/MAINSADR/adrdec2/dec4_3/n8285 , 
        \SADR/MAINSADR/adrdec2/dec4_3/n8287 , 
        \SADR/MAINSADR/adrdec2/dec4_3/n8286 , 
        \SADR/MAINSADR/adrdec2/dec4_3/n8288 , 
        \SADR/MAINSADR/adrdec2/dec4_4/n8283 , 
        \SADR/MAINSADR/adrdec2/dec4_4/n8282 , 
        \SADR/MAINSADR/adrdec2/dec4_4/n8279 , 
        \SADR/MAINSADR/adrdec2/dec4_4/n8280 , 
        \SADR/MAINSADR/adrdec2/dec4_4/n8281 , 
        \SADR/MAINSADR/adrdec2/dec4_5/n8274 , 
        \SADR/MAINSADR/adrdec2/dec4_5/n8275 , 
        \SADR/MAINSADR/adrdec2/dec4_5/n8277 , 
        \SADR/MAINSADR/adrdec2/dec4_5/n8278 , 
        \SADR/MAINSADR/adrdec2/dec4_5/n8276 , 
        \SADR/MAINSADR/adrdec2/dec3_6/n8273 , 
        \SADR/MAINSADR/adrdec2/dec3_6/n8272 , 
        \SADR/MAINSADR/adrdec2/dec3_6/gg_out , 
        \SADR/MAINSADR/adrdec2/dec3_6/n8271 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6966 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6968 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6967 , 
        \REGF/pbmemff21/pbinc19k_1/inc3_5/gp_out , 
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6965 , 
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6964 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6962 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6963 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6961 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6959 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6958 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6960 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6957 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6956 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6953 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6954 , 
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6955 , 
        \SADR/ADDIDX/add_w_x/add0/c_last , \SADR/ADDIDX/add_w_x/add0/n10626 , 
        \SADR/ADDIDX/add_w_x/add0/n10634 , \SADR/ADDIDX/add_w_x/add0/n10641 , 
        \SADR/ADDIDX/add_w_x/add0/n10653 , \SADR/ADDIDX/add_w_x/add0/n10648 , 
        \SADR/ADDIDX/add_w_x/add0/n10623 , \SADR/ADDIDX/add_w_x/add0/n10625 , 
        \SADR/ADDIDX/add_w_x/add0/gp_out , \SADR/ADDIDX/add_w_x/add0/n10628 , 
        \SADR/ADDIDX/add_w_x/add0/n10646 , \SADR/ADDIDX/add_w_x/add0/n10654 , 
        \SADR/ADDIDX/add_w_x/add0/n10629 , \SADR/ADDIDX/add_w_x/add0/n10632 , 
        \SADR/ADDIDX/add_w_x/add0/n10633 , \SADR/ADDIDX/add_w_x/add0/n10635 , 
        \SADR/ADDIDX/add_w_x/add0/n10640 , \SADR/ADDIDX/add_w_x/add0/n10647 , 
        \SADR/ADDIDX/add_w_x/add0/n10649 , \SADR/ADDIDX/add_w_x/add0/n10627 , 
        \SADR/ADDIDX/add_w_x/add0/n10652 , \SADR/ADDIDX/add_w_x/add0/n10637 , 
        \SADR/ADDIDX/add_w_x/add0/n10642 , \SADR/ADDIDX/add_w_x/add0/n10650 , 
        \SADR/ADDIDX/add_w_x/add0/n10630 , \SADR/ADDIDX/add_w_x/add0/n10639 , 
        \SADR/ADDIDX/add_w_x/add0/n10645 , \SADR/ADDIDX/add_w_x/add0/n10638 , 
        \SADR/ADDIDX/add_w_x/add0/n10624 , \SADR/ADDIDX/add_w_x/add0/n10631 , 
        \SADR/ADDIDX/add_w_x/add0/n10636 , \SADR/ADDIDX/add_w_x/add0/n10643 , 
        \SADR/ADDIDX/add_w_x/add0/n10644 , \SADR/ADDIDX/add_w_x/add0/n10651 , 
        \SADR/ADDIDX/add_w_x/add1/c_last , \SADR/ADDIDX/add_w_x/add1/n10594 , 
        \SADR/ADDIDX/add_w_x/add1/n10608 , \SADR/ADDIDX/add_w_x/add1/n10613 , 
        \SADR/ADDIDX/add_w_x/add1/n10601 , \SADR/ADDIDX/add_w_x/add1/n10606 , 
        \SADR/ADDIDX/add_w_x/add1/n10621 , \SADR/ADDIDX/add_w_x/add1/n10591 , 
        \SADR/ADDIDX/add_w_x/add1/n10592 , \SADR/ADDIDX/add_w_x/add1/n10593 , 
        \SADR/ADDIDX/add_w_x/add1/n10607 , \SADR/ADDIDX/add_w_x/add1/n10614 , 
        \SADR/ADDIDX/add_w_x/add1/n10620 , \SADR/ADDIDX/add_w_x/add1/n10615 , 
        \SADR/ADDIDX/add_w_x/add1/n10595 , \SADR/ADDIDX/add_w_x/add1/n10609 , 
        \SADR/ADDIDX/add_w_x/add1/n10612 , \SADR/ADDIDX/add_w_x/add1/n10597 , 
        \SADR/ADDIDX/add_w_x/add1/n10600 , \SADR/ADDIDX/add_w_x/add1/n10610 , 
        \SADR/ADDIDX/add_w_x/add1/n10598 , \SADR/ADDIDX/add_w_x/add1/n10599 , 
        \SADR/ADDIDX/add_w_x/add1/n10602 , \SADR/ADDIDX/add_w_x/add1/n10619 , 
        \SADR/ADDIDX/add_w_x/add1/n10605 , \SADR/ADDIDX/add_w_x/add1/n10617 , 
        \SADR/ADDIDX/add_w_x/add1/n10622 , \SADR/ADDIDX/add_w_x/add1/n10604 , 
        \SADR/ADDIDX/add_w_x/add1/n10616 , \SADR/ADDIDX/add_w_x/add1/n10596 , 
        \SADR/ADDIDX/add_w_x/add1/n10603 , \SADR/ADDIDX/add_w_x/add1/n10611 , 
        \SADR/ADDIDX/add_w_x/add1/n10618 , \SADR/ADDIDX/add_w_x/add2/c_last , 
        \SADR/ADDIDX/add_w_x/add2/n10563 , \SADR/ADDIDX/add_w_x/add2/n10571 , 
        \SADR/ADDIDX/add_w_x/add2/n10586 , \SADR/ADDIDX/add_w_x/add2/n10578 , 
        \SADR/ADDIDX/add_w_x/add2/n10559 , \SADR/ADDIDX/add_w_x/add2/n10564 , 
        \SADR/ADDIDX/add_w_x/add2/n10581 , \SADR/ADDIDX/add_w_x/add2/n10565 , 
        \SADR/ADDIDX/add_w_x/add2/n10576 , \SADR/ADDIDX/add_w_x/add2/n10588 , 
        \SADR/ADDIDX/add_w_x/add2/n10580 , \SADR/ADDIDX/add_w_x/add2/n10560 , 
        \SADR/ADDIDX/add_w_x/add2/n10570 , \SADR/ADDIDX/add_w_x/add2/n10577 , 
        \SADR/ADDIDX/add_w_x/add2/n10589 , \SADR/ADDIDX/add_w_x/add2/n10579 , 
        \SADR/ADDIDX/add_w_x/add2/n10562 , \SADR/ADDIDX/add_w_x/add2/n10587 , 
        \SADR/ADDIDX/add_w_x/add2/n10569 , \SADR/ADDIDX/add_w_x/add2/n10572 , 
        \SADR/ADDIDX/add_w_x/add2/n10561 , \SADR/ADDIDX/add_w_x/add2/n10566 , 
        \SADR/ADDIDX/add_w_x/add2/n10567 , \SADR/ADDIDX/add_w_x/add2/n10582 , 
        \SADR/ADDIDX/add_w_x/add2/n10585 , \SADR/ADDIDX/add_w_x/add2/n10575 , 
        \SADR/ADDIDX/add_w_x/add2/n10590 , \SADR/ADDIDX/add_w_x/add2/n10568 , 
        \SADR/ADDIDX/add_w_x/add2/n10573 , \SADR/ADDIDX/add_w_x/add2/n10574 , 
        \SADR/ADDIDX/add_w_x/add2/n10583 , \SADR/ADDIDX/add_w_x/add2/n10584 , 
        \SADR/ADDIDX/add_w_x/add3/n10531 , \SADR/ADDIDX/add_w_x/add3/n10538 , 
        \SADR/ADDIDX/add_w_x/add3/n10544 , \SADR/ADDIDX/add_w_x/add3/n10556 , 
        \SADR/ADDIDX/add_w_x/add3/n10536 , \SADR/ADDIDX/add_w_x/add3/n10558 , 
        \SADR/ADDIDX/add_w_x/add3/n10527 , \SADR/ADDIDX/add_w_x/add3/n10529 , 
        \SADR/ADDIDX/add_w_x/add3/n10537 , \SADR/ADDIDX/add_w_x/add3/n10542 , 
        \SADR/ADDIDX/add_w_x/add3/n10543 , \SADR/ADDIDX/add_w_x/add3/n10551 , 
        \SADR/ADDIDX/add_w_x/add3/n10539 , \SADR/ADDIDX/add_w_x/add3/n10550 , 
        \SADR/ADDIDX/add_w_x/add3/n10557 , \SADR/ADDIDX/add_w_x/add3/n10530 , 
        \SADR/ADDIDX/add_w_x/add3/n10545 , \SADR/ADDIDX/add_w_x/add3/n10547 , 
        \SADR/ADDIDX/add_w_x/add3/n10555 , \SADR/ADDIDX/add_w_x/add3/n10532 , 
        \SADR/ADDIDX/add_w_x/add3/n10535 , \SADR/ADDIDX/add_w_x/add3/n10540 , 
        \SADR/ADDIDX/add_w_x/add3/n10552 , \SADR/ADDIDX/add_w_x/add3/n10528 , 
        \SADR/ADDIDX/add_w_x/add3/n10533 , \SADR/ADDIDX/add_w_x/add3/n10534 , 
        \SADR/ADDIDX/add_w_x/add3/n10541 , \SADR/ADDIDX/add_w_x/add3/n10549 , 
        \SADR/ADDIDX/add_w_x/add3/n10548 , \SADR/ADDIDX/add_w_x/add3/n10553 , 
        \SADR/ADDIDX/add_w_x/add3/n10554 , \SADR/ADDIDX/add_w_x/add3/n10546 , 
        \SADR/ADDIDX/add_x_z/add0/c_last , \SADR/ADDIDX/add_x_z/add0/n10494 , 
        \SADR/ADDIDX/add_x_z/add0/n10523 , \SADR/ADDIDX/add_x_z/add0/n10504 , 
        \SADR/ADDIDX/add_x_z/add0/n10511 , \SADR/ADDIDX/add_x_z/add0/n10516 , 
        \SADR/ADDIDX/add_x_z/add0/n10495 , \SADR/ADDIDX/add_x_z/add0/n10502 , 
        \SADR/ADDIDX/add_x_z/add0/n10503 , \SADR/ADDIDX/add_x_z/add0/n10518 , 
        \SADR/ADDIDX/add_x_z/add0/n10510 , \SADR/ADDIDX/add_x_z/add0/n10524 , 
        \SADR/ADDIDX/add_x_z/add0/n10505 , \SADR/ADDIDX/add_x_z/add0/n10519 , 
        \SADR/ADDIDX/add_x_z/add0/n10525 , \SADR/ADDIDX/add_x_z/add0/n10522 , 
        \SADR/ADDIDX/add_x_z/add0/n10496 , \SADR/ADDIDX/add_x_z/add0/gp_out , 
        \SADR/ADDIDX/add_x_z/add0/n10497 , \SADR/ADDIDX/add_x_z/add0/n10517 , 
        \SADR/ADDIDX/add_x_z/add0/n10507 , \SADR/ADDIDX/add_x_z/add0/n10498 , 
        \SADR/ADDIDX/add_x_z/add0/n10499 , \SADR/ADDIDX/add_x_z/add0/n10509 , 
        \SADR/ADDIDX/add_x_z/add0/n10512 , \SADR/ADDIDX/add_x_z/add0/n10515 , 
        \SADR/ADDIDX/add_x_z/add0/n10520 , \SADR/ADDIDX/add_x_z/add0/n10500 , 
        \SADR/ADDIDX/add_x_z/add0/n10501 , \SADR/ADDIDX/add_x_z/add0/n10508 , 
        \SADR/ADDIDX/add_x_z/add0/n10513 , \SADR/ADDIDX/add_x_z/add0/n10506 , 
        \SADR/ADDIDX/add_x_z/add0/n10514 , \SADR/ADDIDX/add_x_z/add0/n10521 , 
        \SADR/ADDIDX/add_x_z/add1/c_last , \SADR/ADDIDX/add_x_z/add1/n10471 , 
        \SADR/ADDIDX/add_x_z/add1/n10478 , \SADR/ADDIDX/add_x_z/add1/n10463 , 
        \SADR/ADDIDX/add_x_z/add1/n10486 , \SADR/ADDIDX/add_x_z/add1/n10464 , 
        \SADR/ADDIDX/add_x_z/add1/n10481 , \SADR/ADDIDX/add_x_z/add1/n10462 , 
        \SADR/ADDIDX/add_x_z/add1/n10465 , \SADR/ADDIDX/add_x_z/add1/n10476 , 
        \SADR/ADDIDX/add_x_z/add1/n10488 , \SADR/ADDIDX/add_x_z/add1/n10493 , 
        \SADR/ADDIDX/add_x_z/add1/n10480 , \SADR/ADDIDX/add_x_z/add1/n10470 , 
        \SADR/ADDIDX/add_x_z/add1/n10477 , \SADR/ADDIDX/add_x_z/add1/n10489 , 
        \SADR/ADDIDX/add_x_z/add1/n10492 , \SADR/ADDIDX/add_x_z/add1/n10466 , 
        \SADR/ADDIDX/add_x_z/add1/n10467 , \SADR/ADDIDX/add_x_z/add1/n10479 , 
        \SADR/ADDIDX/add_x_z/add1/n10487 , \SADR/ADDIDX/add_x_z/add1/n10469 , 
        \SADR/ADDIDX/add_x_z/add1/n10472 , \SADR/ADDIDX/add_x_z/add1/n10485 , 
        \SADR/ADDIDX/add_x_z/add1/n10475 , \SADR/ADDIDX/add_x_z/add1/n10482 , 
        \SADR/ADDIDX/add_x_z/add1/n10490 , \SADR/ADDIDX/add_x_z/add1/n10483 , 
        \SADR/ADDIDX/add_x_z/add1/n10468 , \SADR/ADDIDX/add_x_z/add1/n10474 , 
        \SADR/ADDIDX/add_x_z/add1/n10491 , \SADR/ADDIDX/add_x_z/add1/n10473 , 
        \SADR/ADDIDX/add_x_z/add1/n10484 , \SADR/ADDIDX/add_x_z/add2/c_last , 
        \SADR/ADDIDX/add_x_z/add2/n10431 , \SADR/ADDIDX/add_x_z/add2/n10438 , 
        \SADR/ADDIDX/add_x_z/add2/n10456 , \SADR/ADDIDX/add_x_z/add2/n10443 , 
        \SADR/ADDIDX/add_x_z/add2/n10444 , \SADR/ADDIDX/add_x_z/add2/n10430 , 
        \SADR/ADDIDX/add_x_z/add2/n10436 , \SADR/ADDIDX/add_x_z/add2/n10437 , 
        \SADR/ADDIDX/add_x_z/add2/n10451 , \SADR/ADDIDX/add_x_z/add2/n10458 , 
        \SADR/ADDIDX/add_x_z/add2/n10459 , \SADR/ADDIDX/add_x_z/add2/n10439 , 
        \SADR/ADDIDX/add_x_z/add2/n10442 , \SADR/ADDIDX/add_x_z/add2/n10450 , 
        \SADR/ADDIDX/add_x_z/add2/n10445 , \SADR/ADDIDX/add_x_z/add2/n10457 , 
        \SADR/ADDIDX/add_x_z/add2/n10432 , \SADR/ADDIDX/add_x_z/add2/n10455 , 
        \SADR/ADDIDX/add_x_z/add2/n10433 , \SADR/ADDIDX/add_x_z/add2/n10434 , 
        \SADR/ADDIDX/add_x_z/add2/n10435 , \SADR/ADDIDX/add_x_z/add2/n10440 , 
        \SADR/ADDIDX/add_x_z/add2/n10447 , \SADR/ADDIDX/add_x_z/add2/n10460 , 
        \SADR/ADDIDX/add_x_z/add2/n10449 , \SADR/ADDIDX/add_x_z/add2/n10452 , 
        \SADR/ADDIDX/add_x_z/add2/n10441 , \SADR/ADDIDX/add_x_z/add2/n10446 , 
        \SADR/ADDIDX/add_x_z/add2/n10448 , \SADR/ADDIDX/add_x_z/add2/n10453 , 
        \SADR/ADDIDX/add_x_z/add2/n10454 , \SADR/ADDIDX/add_x_z/add2/n10461 , 
        \SADR/ADDIDX/add_x_z/add3/n10404 , \SADR/ADDIDX/add_x_z/add3/n10416 , 
        \SADR/ADDIDX/add_x_z/add3/n10423 , \SADR/ADDIDX/add_x_z/add3/n10398 , 
        \SADR/ADDIDX/add_x_z/add3/n10399 , \SADR/ADDIDX/add_x_z/add3/n10403 , 
        \SADR/ADDIDX/add_x_z/add3/n10411 , \SADR/ADDIDX/add_x_z/add3/n10424 , 
        \SADR/ADDIDX/add_x_z/add3/n10418 , \SADR/ADDIDX/add_x_z/add3/n10410 , 
        \SADR/ADDIDX/add_x_z/add3/n10400 , \SADR/ADDIDX/add_x_z/add3/n10402 , 
        \SADR/ADDIDX/add_x_z/add3/n10419 , \SADR/ADDIDX/add_x_z/add3/n10425 , 
        \SADR/ADDIDX/add_x_z/add3/n10405 , \SADR/ADDIDX/add_x_z/add3/n10422 , 
        \SADR/ADDIDX/add_x_z/add3/n10417 , \SADR/ADDIDX/add_x_z/add3/n10407 , 
        \SADR/ADDIDX/add_x_z/add3/n10420 , \SADR/ADDIDX/add_x_z/add3/n10409 , 
        \SADR/ADDIDX/add_x_z/add3/n10415 , \SADR/ADDIDX/add_x_z/add3/n10429 , 
        \SADR/ADDIDX/add_x_z/add3/n10412 , \SADR/ADDIDX/add_x_z/add3/n10401 , 
        \SADR/ADDIDX/add_x_z/add3/n10408 , \SADR/ADDIDX/add_x_z/add3/n10413 , 
        \SADR/ADDIDX/add_x_z/add3/n10427 , \SADR/ADDIDX/add_x_z/add3/n10406 , 
        \SADR/ADDIDX/add_x_z/add3/n10421 , \SADR/ADDIDX/add_x_z/add3/n10426 , 
        \SADR/ADDIDX/add_x_z/add3/n10414 , \SADR/ADDIDX/add_x_z/add3/n10428 , 
        \SADR/ADDIDX/add_y_z/add0/c_last , \SADR/ADDIDX/add_y_z/add0/n10372 , 
        \SADR/ADDIDX/add_y_z/add0/n10385 , \SADR/ADDIDX/add_y_z/add0/n10369 , 
        \SADR/ADDIDX/add_y_z/add0/n10365 , \SADR/ADDIDX/add_y_z/add0/n10366 , 
        \SADR/ADDIDX/add_y_z/add0/n10367 , \SADR/ADDIDX/add_y_z/add0/n10375 , 
        \SADR/ADDIDX/add_y_z/add0/n10390 , \SADR/ADDIDX/add_y_z/add0/n10374 , 
        \SADR/ADDIDX/add_y_z/add0/n10382 , \SADR/ADDIDX/add_y_z/add0/n10383 , 
        \SADR/ADDIDX/add_y_z/add0/n10391 , \SADR/ADDIDX/add_y_z/add0/gp_out , 
        \SADR/ADDIDX/add_y_z/add0/n10368 , \SADR/ADDIDX/add_y_z/add0/n10384 , 
        \SADR/ADDIDX/add_y_z/add0/n10371 , \SADR/ADDIDX/add_y_z/add0/n10373 , 
        \SADR/ADDIDX/add_y_z/add0/n10396 , \SADR/ADDIDX/add_y_z/add0/n10378 , 
        \SADR/ADDIDX/add_y_z/add0/n10386 , \SADR/ADDIDX/add_y_z/add0/n10376 , 
        \SADR/ADDIDX/add_y_z/add0/n10388 , \SADR/ADDIDX/add_y_z/add0/n10394 , 
        \SADR/ADDIDX/add_y_z/add0/n10393 , \SADR/ADDIDX/add_y_z/add0/n10377 , 
        \SADR/ADDIDX/add_y_z/add0/n10381 , \SADR/ADDIDX/add_y_z/add0/n10380 , 
        \SADR/ADDIDX/add_y_z/add0/n10389 , \SADR/ADDIDX/add_y_z/add0/n10392 , 
        \SADR/ADDIDX/add_y_z/add0/n10370 , \SADR/ADDIDX/add_y_z/add0/n10379 , 
        \SADR/ADDIDX/add_y_z/add0/n10387 , \SADR/ADDIDX/add_y_z/add0/n10395 , 
        \SADR/ADDIDX/add_y_z/add1/c_last , \SADR/ADDIDX/add_y_z/add1/n10347 , 
        \SADR/ADDIDX/add_y_z/add1/n10355 , \SADR/ADDIDX/add_y_z/add1/n10360 , 
        \SADR/ADDIDX/add_y_z/add1/n10349 , \SADR/ADDIDX/add_y_z/add1/n10333 , 
        \SADR/ADDIDX/add_y_z/add1/n10334 , \SADR/ADDIDX/add_y_z/add1/n10335 , 
        \SADR/ADDIDX/add_y_z/add1/n10340 , \SADR/ADDIDX/add_y_z/add1/n10352 , 
        \SADR/ADDIDX/add_y_z/add1/n10348 , \SADR/ADDIDX/add_y_z/add1/n10353 , 
        \SADR/ADDIDX/add_y_z/add1/n10341 , \SADR/ADDIDX/add_y_z/add1/n10346 , 
        \SADR/ADDIDX/add_y_z/add1/n10361 , \SADR/ADDIDX/add_y_z/add1/n10336 , 
        \SADR/ADDIDX/add_y_z/add1/n10338 , \SADR/ADDIDX/add_y_z/add1/n10354 , 
        \SADR/ADDIDX/add_y_z/add1/n10344 , \SADR/ADDIDX/add_y_z/add1/n10363 , 
        \SADR/ADDIDX/add_y_z/add1/n10356 , \SADR/ADDIDX/add_y_z/add1/n10343 , 
        \SADR/ADDIDX/add_y_z/add1/n10351 , \SADR/ADDIDX/add_y_z/add1/n10364 , 
        \SADR/ADDIDX/add_y_z/add1/n10337 , \SADR/ADDIDX/add_y_z/add1/n10350 , 
        \SADR/ADDIDX/add_y_z/add1/n10358 , \SADR/ADDIDX/add_y_z/add1/n10359 , 
        \SADR/ADDIDX/add_y_z/add1/n10339 , \SADR/ADDIDX/add_y_z/add1/n10342 , 
        \SADR/ADDIDX/add_y_z/add1/n10345 , \SADR/ADDIDX/add_y_z/add1/n10362 , 
        \SADR/ADDIDX/add_y_z/add1/n10357 , \SADR/ADDIDX/add_y_z/add2/c_last , 
        \SADR/ADDIDX/add_y_z/add2/n10315 , \SADR/ADDIDX/add_y_z/add2/n10332 , 
        \SADR/ADDIDX/add_y_z/add2/n10320 , \SADR/ADDIDX/add_y_z/add2/n10329 , 
        \SADR/ADDIDX/add_y_z/add2/n10307 , \SADR/ADDIDX/add_y_z/add2/n10327 , 
        \SADR/ADDIDX/add_y_z/add2/n10301 , \SADR/ADDIDX/add_y_z/add2/n10309 , 
        \SADR/ADDIDX/add_y_z/add2/n10312 , \SADR/ADDIDX/add_y_z/add2/n10302 , 
        \SADR/ADDIDX/add_y_z/add2/n10303 , \SADR/ADDIDX/add_y_z/add2/n10308 , 
        \SADR/ADDIDX/add_y_z/add2/n10313 , \SADR/ADDIDX/add_y_z/add2/n10326 , 
        \SADR/ADDIDX/add_y_z/add2/n10314 , \SADR/ADDIDX/add_y_z/add2/n10328 , 
        \SADR/ADDIDX/add_y_z/add2/n10304 , \SADR/ADDIDX/add_y_z/add2/n10306 , 
        \SADR/ADDIDX/add_y_z/add2/n10321 , \SADR/ADDIDX/add_y_z/add2/n10316 , 
        \SADR/ADDIDX/add_y_z/add2/n10331 , \SADR/ADDIDX/add_y_z/add2/n10323 , 
        \SADR/ADDIDX/add_y_z/add2/n10324 , \SADR/ADDIDX/add_y_z/add2/n10311 , 
        \SADR/ADDIDX/add_y_z/add2/n10318 , \SADR/ADDIDX/add_y_z/add2/n10319 , 
        \SADR/ADDIDX/add_y_z/add2/n10325 , \SADR/ADDIDX/add_y_z/add2/n10305 , 
        \SADR/ADDIDX/add_y_z/add2/n10310 , \SADR/ADDIDX/add_y_z/add2/n10317 , 
        \SADR/ADDIDX/add_y_z/add2/n10330 , \SADR/ADDIDX/add_y_z/add2/n10322 , 
        \SADR/ADDIDX/add_y_z/add3/n10269 , \SADR/ADDIDX/add_y_z/add3/n10285 , 
        \SADR/ADDIDX/add_y_z/add3/n10272 , \SADR/ADDIDX/add_y_z/add3/n10297 , 
        \SADR/ADDIDX/add_y_z/add3/n10275 , \SADR/ADDIDX/add_y_z/add3/n10290 , 
        \SADR/ADDIDX/add_y_z/add3/n10300 , \SADR/ADDIDX/add_y_z/add3/n10270 , 
        \SADR/ADDIDX/add_y_z/add3/n10271 , \SADR/ADDIDX/add_y_z/add3/n10273 , 
        \SADR/ADDIDX/add_y_z/add3/n10274 , \SADR/ADDIDX/add_y_z/add3/n10282 , 
        \SADR/ADDIDX/add_y_z/add3/n10299 , \SADR/ADDIDX/add_y_z/add3/n10291 , 
        \SADR/ADDIDX/add_y_z/add3/n10283 , \SADR/ADDIDX/add_y_z/add3/n10284 , 
        \SADR/ADDIDX/add_y_z/add3/n10298 , \SADR/ADDIDX/add_y_z/add3/n10296 , 
        \SADR/ADDIDX/add_y_z/add3/n10278 , \SADR/ADDIDX/add_y_z/add3/n10286 , 
        \SADR/ADDIDX/add_y_z/add3/n10294 , \SADR/ADDIDX/add_y_z/add3/n10276 , 
        \SADR/ADDIDX/add_y_z/add3/n10277 , \SADR/ADDIDX/add_y_z/add3/n10281 , 
        \SADR/ADDIDX/add_y_z/add3/n10288 , \SADR/ADDIDX/add_y_z/add3/n10293 , 
        \SADR/ADDIDX/add_y_z/add3/n10289 , \SADR/ADDIDX/add_y_z/add3/n10292 , 
        \SADR/ADDIDX/add_y_z/add3/n10279 , \SADR/ADDIDX/add_y_z/add3/n10280 , 
        \SADR/ADDIDX/add_y_z/add3/n10287 , \SADR/ADDIDX/add_y_z/add3/n10295 , 
        \SADR/ADDIDX/add_w_y/add0/c_last , \SADR/ADDIDX/add_w_y/add0/n10247 , 
        \SADR/ADDIDX/add_w_y/add0/n10260 , \SADR/ADDIDX/add_w_y/add0/n10252 , 
        \SADR/ADDIDX/add_w_y/add0/n10255 , \SADR/ADDIDX/add_w_y/add0/n10236 , 
        \SADR/ADDIDX/add_w_y/add0/n10238 , \SADR/ADDIDX/add_w_y/add0/gp_out , 
        \SADR/ADDIDX/add_w_y/add0/n10240 , \SADR/ADDIDX/add_w_y/add0/n10249 , 
        \SADR/ADDIDX/add_w_y/add0/n10241 , \SADR/ADDIDX/add_w_y/add0/n10248 , 
        \SADR/ADDIDX/add_w_y/add0/n10267 , \SADR/ADDIDX/add_w_y/add0/n10253 , 
        \SADR/ADDIDX/add_w_y/add0/n10246 , \SADR/ADDIDX/add_w_y/add0/n10266 , 
        \SADR/ADDIDX/add_w_y/add0/n10261 , \SADR/ADDIDX/add_w_y/add0/n10254 , 
        \SADR/ADDIDX/add_w_y/add0/n10244 , \SADR/ADDIDX/add_w_y/add0/n10263 , 
        \SADR/ADDIDX/add_w_y/add0/n10251 , \SADR/ADDIDX/add_w_y/add0/n10256 , 
        \SADR/ADDIDX/add_w_y/add0/n10258 , \SADR/ADDIDX/add_w_y/add0/n10237 , 
        \SADR/ADDIDX/add_w_y/add0/n10242 , \SADR/ADDIDX/add_w_y/add0/n10243 , 
        \SADR/ADDIDX/add_w_y/add0/n10264 , \SADR/ADDIDX/add_w_y/add0/n10250 , 
        \SADR/ADDIDX/add_w_y/add0/n10265 , \SADR/ADDIDX/add_w_y/add0/n10239 , 
        \SADR/ADDIDX/add_w_y/add0/n10245 , \SADR/ADDIDX/add_w_y/add0/n10259 , 
        \SADR/ADDIDX/add_w_y/add0/n10257 , \SADR/ADDIDX/add_w_y/add0/n10262 , 
        \SADR/ADDIDX/add_w_y/add1/c_last , \SADR/ADDIDX/add_w_y/add1/n10207 , 
        \SADR/ADDIDX/add_w_y/add1/n10215 , \SADR/ADDIDX/add_w_y/add1/n10229 , 
        \SADR/ADDIDX/add_w_y/add1/n10232 , \SADR/ADDIDX/add_w_y/add1/n10220 , 
        \SADR/ADDIDX/add_w_y/add1/n10204 , \SADR/ADDIDX/add_w_y/add1/n10206 , 
        \SADR/ADDIDX/add_w_y/add1/n10208 , \SADR/ADDIDX/add_w_y/add1/n10209 , 
        \SADR/ADDIDX/add_w_y/add1/n10212 , \SADR/ADDIDX/add_w_y/add1/n10227 , 
        \SADR/ADDIDX/add_w_y/add1/n10235 , \SADR/ADDIDX/add_w_y/add1/n10226 , 
        \SADR/ADDIDX/add_w_y/add1/n10213 , \SADR/ADDIDX/add_w_y/add1/n10234 , 
        \SADR/ADDIDX/add_w_y/add1/n10214 , \SADR/ADDIDX/add_w_y/add1/n10228 , 
        \SADR/ADDIDX/add_w_y/add1/n10233 , \SADR/ADDIDX/add_w_y/add1/n10221 , 
        \SADR/ADDIDX/add_w_y/add1/n10216 , \SADR/ADDIDX/add_w_y/add1/n10231 , 
        \SADR/ADDIDX/add_w_y/add1/n10223 , \SADR/ADDIDX/add_w_y/add1/n10205 , 
        \SADR/ADDIDX/add_w_y/add1/n10210 , \SADR/ADDIDX/add_w_y/add1/n10211 , 
        \SADR/ADDIDX/add_w_y/add1/n10218 , \SADR/ADDIDX/add_w_y/add1/n10224 , 
        \SADR/ADDIDX/add_w_y/add1/n10219 , \SADR/ADDIDX/add_w_y/add1/n10225 , 
        \SADR/ADDIDX/add_w_y/add1/n10217 , \SADR/ADDIDX/add_w_y/add1/n10230 , 
        \SADR/ADDIDX/add_w_y/add1/n10222 , \SADR/ADDIDX/add_w_y/add2/c_last , 
        \SADR/ADDIDX/add_w_y/add2/n10177 , \SADR/ADDIDX/add_w_y/add2/n10180 , 
        \SADR/ADDIDX/add_w_y/add2/n10189 , \SADR/ADDIDX/add_w_y/add2/n10192 , 
        \SADR/ADDIDX/add_w_y/add2/n10187 , \SADR/ADDIDX/add_w_y/add2/n10172 , 
        \SADR/ADDIDX/add_w_y/add2/n10173 , \SADR/ADDIDX/add_w_y/add2/n10174 , 
        \SADR/ADDIDX/add_w_y/add2/n10176 , \SADR/ADDIDX/add_w_y/add2/n10178 , 
        \SADR/ADDIDX/add_w_y/add2/n10179 , \SADR/ADDIDX/add_w_y/add2/n10200 , 
        \SADR/ADDIDX/add_w_y/add2/n10195 , \SADR/ADDIDX/add_w_y/add2/n10186 , 
        \SADR/ADDIDX/add_w_y/add2/n10201 , \SADR/ADDIDX/add_w_y/add2/n10188 , 
        \SADR/ADDIDX/add_w_y/add2/n10194 , \SADR/ADDIDX/add_w_y/add2/n10193 , 
        \SADR/ADDIDX/add_w_y/add2/n10181 , \SADR/ADDIDX/add_w_y/add2/n10183 , 
        \SADR/ADDIDX/add_w_y/add2/n10191 , \SADR/ADDIDX/add_w_y/add2/n10198 , 
        \SADR/ADDIDX/add_w_y/add2/n10184 , \SADR/ADDIDX/add_w_y/add2/n10196 , 
        \SADR/ADDIDX/add_w_y/add2/n10203 , \SADR/ADDIDX/add_w_y/add2/n10185 , 
        \SADR/ADDIDX/add_w_y/add2/n10202 , \SADR/ADDIDX/add_w_y/add2/n10175 , 
        \SADR/ADDIDX/add_w_y/add2/n10190 , \SADR/ADDIDX/add_w_y/add2/n10197 , 
        \SADR/ADDIDX/add_w_y/add2/n10182 , \SADR/ADDIDX/add_w_y/add2/n10199 , 
        \SADR/ADDIDX/add_w_y/add3/n10150 , \SADR/ADDIDX/add_w_y/add3/n10159 , 
        \SADR/ADDIDX/add_w_y/add3/n10142 , \SADR/ADDIDX/add_w_y/add3/n10145 , 
        \SADR/ADDIDX/add_w_y/add3/n10162 , \SADR/ADDIDX/add_w_y/add3/n10165 , 
        \SADR/ADDIDX/add_w_y/add3/n10140 , \SADR/ADDIDX/add_w_y/add3/n10141 , 
        \SADR/ADDIDX/add_w_y/add3/n10143 , \SADR/ADDIDX/add_w_y/add3/n10144 , 
        \SADR/ADDIDX/add_w_y/add3/n10157 , \SADR/ADDIDX/add_w_y/add3/n10170 , 
        \SADR/ADDIDX/add_w_y/add3/n10163 , \SADR/ADDIDX/add_w_y/add3/n10151 , 
        \SADR/ADDIDX/add_w_y/add3/n10156 , \SADR/ADDIDX/add_w_y/add3/n10171 , 
        \SADR/ADDIDX/add_w_y/add3/n10164 , \SADR/ADDIDX/add_w_y/add3/n10148 , 
        \SADR/ADDIDX/add_w_y/add3/n10153 , \SADR/ADDIDX/add_w_y/add3/n10158 , 
        \SADR/ADDIDX/add_w_y/add3/n10166 , \SADR/ADDIDX/add_w_y/add3/n10146 , 
        \SADR/ADDIDX/add_w_y/add3/n10147 , \SADR/ADDIDX/add_w_y/add3/n10154 , 
        \SADR/ADDIDX/add_w_y/add3/n10161 , \SADR/ADDIDX/add_w_y/add3/n10168 , 
        \SADR/ADDIDX/add_w_y/add3/n10149 , \SADR/ADDIDX/add_w_y/add3/n10155 , 
        \SADR/ADDIDX/add_w_y/add3/n10160 , \SADR/ADDIDX/add_w_y/add3/n10169 , 
        \SADR/ADDIDX/add_w_y/add3/n10152 , \SADR/ADDIDX/add_w_y/add3/n10167 , 
        \SADR/ADDIDX/add_w_x_y/add0/c_last , 
        \SADR/ADDIDX/add_w_x_y/add0/n10110 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10119 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10125 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10137 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10107 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10108 , 
        \SADR/ADDIDX/add_w_x_y/add0/gp_out , 
        \SADR/ADDIDX/add_w_x_y/add0/n10116 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10117 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10122 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10130 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10118 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10123 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10131 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10138 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10124 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10111 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10136 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10113 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10126 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10134 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10114 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10128 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10133 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10115 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10121 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10132 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10120 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10129 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10109 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10127 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10112 , 
        \SADR/ADDIDX/add_w_x_y/add0/n10135 , 
        \SADR/ADDIDX/add_w_x_y/add1/c_last , 
        \SADR/ADDIDX/add_w_x_y/add1/n10077 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10089 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10092 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10102 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10080 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10079 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10075 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10076 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10078 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10086 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10087 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10095 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10105 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10094 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10104 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10088 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10093 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10103 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10081 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10083 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10091 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10101 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10084 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10098 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10085 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10096 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10106 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10097 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10082 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10090 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10100 , 
        \SADR/ADDIDX/add_w_x_y/add1/n10099 , 
        \SADR/ADDIDX/add_w_x_y/add2/c_last , 
        \SADR/ADDIDX/add_w_x_y/add2/n10050 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10065 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10059 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10043 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10044 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10045 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10057 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10062 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10070 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10051 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10056 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10063 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10071 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10058 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10064 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10046 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10048 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10053 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10061 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10074 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10066 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10047 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10054 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10073 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10060 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10068 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10049 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10052 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10055 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10069 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10072 , 
        \SADR/ADDIDX/add_w_x_y/add2/n10067 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10019 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10025 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10037 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10042 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10017 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10030 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10011 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10016 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10022 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10039 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10031 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10018 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10023 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10038 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10024 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10012 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10013 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10036 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10026 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10034 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10041 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10014 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10015 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10021 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10028 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10033 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10029 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10020 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10032 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10027 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10035 , 
        \SADR/ADDIDX/add_w_x_y/add3/n10040 , 
        \SADR/ADDIDX/add_x_y_z/add0/c_last , 
        \SADR/ADDIDX/add_x_y_z/add0/n9978 , \SADR/ADDIDX/add_x_y_z/add0/n9986 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10002 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9994 , \SADR/ADDIDX/add_x_y_z/add0/n9988 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9979 , \SADR/ADDIDX/add_x_y_z/add0/n9980 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9981 , \SADR/ADDIDX/add_x_y_z/add0/n9993 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9989 , \SADR/ADDIDX/add_x_y_z/add0/n9992 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10005 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10004 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9987 , 
        \SADR/ADDIDX/add_x_y_z/add0/gp_out , 
        \SADR/ADDIDX/add_x_y_z/add0/n10003 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9982 , \SADR/ADDIDX/add_x_y_z/add0/n9995 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9985 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10001 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9990 , \SADR/ADDIDX/add_x_y_z/add0/n9997 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10008 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9983 , \SADR/ADDIDX/add_x_y_z/add0/n9991 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9999 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10006 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9998 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10007 , 
        \SADR/ADDIDX/add_x_y_z/add0/n9984 , \SADR/ADDIDX/add_x_y_z/add0/n9996 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10000 , 
        \SADR/ADDIDX/add_x_y_z/add0/n10009 , 
        \SADR/ADDIDX/add_x_y_z/add1/c_last , 
        \SADR/ADDIDX/add_x_y_z/add1/n9956 , \SADR/ADDIDX/add_x_y_z/add1/n9963 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9971 , \SADR/ADDIDX/add_x_y_z/add1/n9946 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9947 , \SADR/ADDIDX/add_x_y_z/add1/n9950 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9951 , \SADR/ADDIDX/add_x_y_z/add1/n9958 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9964 , \SADR/ADDIDX/add_x_y_z/add1/n9976 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9959 , \SADR/ADDIDX/add_x_y_z/add1/n9977 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9962 , \SADR/ADDIDX/add_x_y_z/add1/n9965 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9957 , \SADR/ADDIDX/add_x_y_z/add1/n9970 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9948 , \SADR/ADDIDX/add_x_y_z/add1/n9949 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9955 , \SADR/ADDIDX/add_x_y_z/add1/n9960 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9969 , \SADR/ADDIDX/add_x_y_z/add1/n9972 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9952 , \SADR/ADDIDX/add_x_y_z/add1/n9975 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9953 , \SADR/ADDIDX/add_x_y_z/add1/n9967 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9974 , \SADR/ADDIDX/add_x_y_z/add1/n9966 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9954 , \SADR/ADDIDX/add_x_y_z/add1/n9961 , 
        \SADR/ADDIDX/add_x_y_z/add1/n9968 , \SADR/ADDIDX/add_x_y_z/add1/n9973 , 
        \SADR/ADDIDX/add_x_y_z/add2/c_last , 
        \SADR/ADDIDX/add_x_y_z/add2/n9916 , \SADR/ADDIDX/add_x_y_z/add2/n9931 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9938 , \SADR/ADDIDX/add_x_y_z/add2/n9944 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9923 , \SADR/ADDIDX/add_x_y_z/add2/n9924 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9914 , \SADR/ADDIDX/add_x_y_z/add2/n9915 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9917 , \SADR/ADDIDX/add_x_y_z/add2/n9918 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9919 , \SADR/ADDIDX/add_x_y_z/add2/n9936 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9943 , \SADR/ADDIDX/add_x_y_z/add2/n9925 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9937 , \SADR/ADDIDX/add_x_y_z/add2/n9942 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9945 , \SADR/ADDIDX/add_x_y_z/add2/n9922 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9930 , \SADR/ADDIDX/add_x_y_z/add2/n9939 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9932 , \SADR/ADDIDX/add_x_y_z/add2/n9920 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9929 , \SADR/ADDIDX/add_x_y_z/add2/n9926 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9927 , \SADR/ADDIDX/add_x_y_z/add2/n9935 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9940 , \SADR/ADDIDX/add_x_y_z/add2/n9928 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9934 , \SADR/ADDIDX/add_x_y_z/add2/n9941 , 
        \SADR/ADDIDX/add_x_y_z/add2/n9933 , \SADR/ADDIDX/add_x_y_z/add2/n9921 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9886 , \SADR/ADDIDX/add_x_y_z/add3/n9893 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9894 , \SADR/ADDIDX/add_x_y_z/add3/n9904 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9903 , \SADR/ADDIDX/add_x_y_z/add3/n9882 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9887 , \SADR/ADDIDX/add_x_y_z/add3/n9888 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9889 , \SADR/ADDIDX/add_x_y_z/add3/n9911 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9892 , \SADR/ADDIDX/add_x_y_z/add3/n9902 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9910 , \SADR/ADDIDX/add_x_y_z/add3/n9895 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9905 , \SADR/ADDIDX/add_x_y_z/add3/n9885 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9890 , \SADR/ADDIDX/add_x_y_z/add3/n9897 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9900 , \SADR/ADDIDX/add_x_y_z/add3/n9907 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9899 , \SADR/ADDIDX/add_x_y_z/add3/n9909 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9883 , \SADR/ADDIDX/add_x_y_z/add3/n9891 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9912 , \SADR/ADDIDX/add_x_y_z/add3/n9901 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9913 , \SADR/ADDIDX/add_x_y_z/add3/n9884 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9898 , \SADR/ADDIDX/add_x_y_z/add3/n9908 , 
        \SADR/ADDIDX/add_x_y_z/add3/n9896 , \SADR/ADDIDX/add_x_y_z/add3/n9906 , 
        \SADR/ADDIDX/add_w_z/add0/c_last , \SADR/ADDIDX/add_w_z/add0/n9856 , 
        \SADR/ADDIDX/add_w_z/add0/n9863 , \SADR/ADDIDX/add_w_z/add0/n9878 , 
        \SADR/ADDIDX/add_w_z/add0/n9871 , \SADR/ADDIDX/add_w_z/add0/n9851 , 
        \SADR/ADDIDX/add_w_z/add0/n9876 , \SADR/ADDIDX/add_w_z/add0/n9849 , 
        \SADR/ADDIDX/add_w_z/add0/n9850 , \SADR/ADDIDX/add_w_z/add0/n9858 , 
        \SADR/ADDIDX/add_w_z/add0/n9864 , \SADR/ADDIDX/add_w_z/add0/n9877 , 
        \SADR/ADDIDX/add_w_z/add0/gp_out , \SADR/ADDIDX/add_w_z/add0/n9859 , 
        \SADR/ADDIDX/add_w_z/add0/n9865 , \SADR/ADDIDX/add_w_z/add0/n9880 , 
        \SADR/ADDIDX/add_w_z/add0/n9862 , \SADR/ADDIDX/add_w_z/add0/n9879 , 
        \SADR/ADDIDX/add_w_z/add0/n9852 , \SADR/ADDIDX/add_w_z/add0/n9855 , 
        \SADR/ADDIDX/add_w_z/add0/n9857 , \SADR/ADDIDX/add_w_z/add0/n9870 , 
        \SADR/ADDIDX/add_w_z/add0/n9860 , \SADR/ADDIDX/add_w_z/add0/n9869 , 
        \SADR/ADDIDX/add_w_z/add0/n9872 , \SADR/ADDIDX/add_w_z/add0/n9875 , 
        \SADR/ADDIDX/add_w_z/add0/n9853 , \SADR/ADDIDX/add_w_z/add0/n9867 , 
        \SADR/ADDIDX/add_w_z/add0/n9854 , \SADR/ADDIDX/add_w_z/add0/n9861 , 
        \SADR/ADDIDX/add_w_z/add0/n9866 , \SADR/ADDIDX/add_w_z/add0/n9874 , 
        \SADR/ADDIDX/add_w_z/add0/n9873 , \SADR/ADDIDX/add_w_z/add0/n9868 , 
        \SADR/ADDIDX/add_w_z/add1/c_last , \SADR/ADDIDX/add_w_z/add1/n9823 , 
        \SADR/ADDIDX/add_w_z/add1/n9831 , \SADR/ADDIDX/add_w_z/add1/n9844 , 
        \SADR/ADDIDX/add_w_z/add1/n9818 , \SADR/ADDIDX/add_w_z/add1/n9838 , 
        \SADR/ADDIDX/add_w_z/add1/n9817 , \SADR/ADDIDX/add_w_z/add1/n9819 , 
        \SADR/ADDIDX/add_w_z/add1/n9824 , \SADR/ADDIDX/add_w_z/add1/n9825 , 
        \SADR/ADDIDX/add_w_z/add1/n9836 , \SADR/ADDIDX/add_w_z/add1/n9843 , 
        \SADR/ADDIDX/add_w_z/add1/n9830 , \SADR/ADDIDX/add_w_z/add1/n9837 , 
        \SADR/ADDIDX/add_w_z/add1/n9842 , \SADR/ADDIDX/add_w_z/add1/n9845 , 
        \SADR/ADDIDX/add_w_z/add1/n9820 , \SADR/ADDIDX/add_w_z/add1/n9822 , 
        \SADR/ADDIDX/add_w_z/add1/n9839 , \SADR/ADDIDX/add_w_z/add1/n9829 , 
        \SADR/ADDIDX/add_w_z/add1/n9832 , \SADR/ADDIDX/add_w_z/add1/n9847 , 
        \SADR/ADDIDX/add_w_z/add1/n9821 , \SADR/ADDIDX/add_w_z/add1/n9826 , 
        \SADR/ADDIDX/add_w_z/add1/n9827 , \SADR/ADDIDX/add_w_z/add1/n9835 , 
        \SADR/ADDIDX/add_w_z/add1/n9840 , \SADR/ADDIDX/add_w_z/add1/n9828 , 
        \SADR/ADDIDX/add_w_z/add1/n9833 , \SADR/ADDIDX/add_w_z/add1/n9834 , 
        \SADR/ADDIDX/add_w_z/add1/n9841 , \SADR/ADDIDX/add_w_z/add1/n9848 , 
        \SADR/ADDIDX/add_w_z/add1/n9846 , \SADR/ADDIDX/add_w_z/add2/c_last , 
        \SADR/ADDIDX/add_w_z/add2/n9796 , \SADR/ADDIDX/add_w_z/add2/n9804 , 
        \SADR/ADDIDX/add_w_z/add2/n9816 , \SADR/ADDIDX/add_w_z/add2/n9785 , 
        \SADR/ADDIDX/add_w_z/add2/n9790 , \SADR/ADDIDX/add_w_z/add2/n9791 , 
        \SADR/ADDIDX/add_w_z/add2/n9798 , \SADR/ADDIDX/add_w_z/add2/n9803 , 
        \SADR/ADDIDX/add_w_z/add2/n9811 , \SADR/ADDIDX/add_w_z/add2/n9799 , 
        \SADR/ADDIDX/add_w_z/add2/n9802 , \SADR/ADDIDX/add_w_z/add2/n9797 , 
        \SADR/ADDIDX/add_w_z/add2/n9810 , \SADR/ADDIDX/add_w_z/add2/n9786 , 
        \SADR/ADDIDX/add_w_z/add2/n9787 , \SADR/ADDIDX/add_w_z/add2/n9805 , 
        \SADR/ADDIDX/add_w_z/add2/n9795 , \SADR/ADDIDX/add_w_z/add2/n9815 , 
        \SADR/ADDIDX/add_w_z/add2/n9807 , \SADR/ADDIDX/add_w_z/add2/n9788 , 
        \SADR/ADDIDX/add_w_z/add2/n9789 , \SADR/ADDIDX/add_w_z/add2/n9792 , 
        \SADR/ADDIDX/add_w_z/add2/n9800 , \SADR/ADDIDX/add_w_z/add2/n9812 , 
        \SADR/ADDIDX/add_w_z/add2/n9801 , \SADR/ADDIDX/add_w_z/add2/n9809 , 
        \SADR/ADDIDX/add_w_z/add2/n9808 , \SADR/ADDIDX/add_w_z/add2/n9793 , 
        \SADR/ADDIDX/add_w_z/add2/n9794 , \SADR/ADDIDX/add_w_z/add2/n9813 , 
        \SADR/ADDIDX/add_w_z/add2/n9814 , \SADR/ADDIDX/add_w_z/add2/n9806 , 
        \SADR/ADDIDX/add_w_z/add3/n9754 , \SADR/ADDIDX/add_w_z/add3/n9768 , 
        \SADR/ADDIDX/add_w_z/add3/n9773 , \SADR/ADDIDX/add_w_z/add3/n9761 , 
        \SADR/ADDIDX/add_w_z/add3/n9784 , \SADR/ADDIDX/add_w_z/add3/n9753 , 
        \SADR/ADDIDX/add_w_z/add3/n9766 , \SADR/ADDIDX/add_w_z/add3/n9783 , 
        \SADR/ADDIDX/add_w_z/add3/n9755 , \SADR/ADDIDX/add_w_z/add3/n9767 , 
        \SADR/ADDIDX/add_w_z/add3/n9774 , \SADR/ADDIDX/add_w_z/add3/n9772 , 
        \SADR/ADDIDX/add_w_z/add3/n9782 , \SADR/ADDIDX/add_w_z/add3/n9775 , 
        \SADR/ADDIDX/add_w_z/add3/n9769 , \SADR/ADDIDX/add_w_z/add3/n9756 , 
        \SADR/ADDIDX/add_w_z/add3/n9757 , \SADR/ADDIDX/add_w_z/add3/n9760 , 
        \SADR/ADDIDX/add_w_z/add3/n9758 , \SADR/ADDIDX/add_w_z/add3/n9759 , 
        \SADR/ADDIDX/add_w_z/add3/n9762 , \SADR/ADDIDX/add_w_z/add3/n9770 , 
        \SADR/ADDIDX/add_w_z/add3/n9779 , \SADR/ADDIDX/add_w_z/add3/n9764 , 
        \SADR/ADDIDX/add_w_z/add3/n9765 , \SADR/ADDIDX/add_w_z/add3/n9780 , 
        \SADR/ADDIDX/add_w_z/add3/n9777 , \SADR/ADDIDX/add_w_z/add3/n9781 , 
        \SADR/ADDIDX/add_w_z/add3/n9776 , \SADR/ADDIDX/add_w_z/add3/n9763 , 
        \SADR/ADDIDX/add_w_z/add3/n9771 , \SADR/ADDIDX/add_w_z/add3/n9778 , 
        \SADR/ADDIDX/add_x_y/add0/c_last , \SADR/ADDIDX/add_x_y/add0/n9721 , 
        \SADR/ADDIDX/add_x_y/add0/n9728 , \SADR/ADDIDX/add_x_y/add0/n9746 , 
        \SADR/ADDIDX/add_x_y/add0/n9733 , \SADR/ADDIDX/add_x_y/add0/n9734 , 
        \SADR/ADDIDX/add_x_y/add0/n9720 , \SADR/ADDIDX/add_x_y/add0/n9726 , 
        \SADR/ADDIDX/add_x_y/add0/n9741 , \SADR/ADDIDX/add_x_y/add0/n9727 , 
        \SADR/ADDIDX/add_x_y/add0/n9735 , \SADR/ADDIDX/add_x_y/add0/n9740 , 
        \SADR/ADDIDX/add_x_y/add0/n9748 , \SADR/ADDIDX/add_x_y/add0/n9749 , 
        \SADR/ADDIDX/add_x_y/add0/n9722 , \SADR/ADDIDX/add_x_y/add0/gp_out , 
        \SADR/ADDIDX/add_x_y/add0/n9729 , \SADR/ADDIDX/add_x_y/add0/n9732 , 
        \SADR/ADDIDX/add_x_y/add0/n9747 , \SADR/ADDIDX/add_x_y/add0/n9723 , 
        \SADR/ADDIDX/add_x_y/add0/n9724 , \SADR/ADDIDX/add_x_y/add0/n9725 , 
        \SADR/ADDIDX/add_x_y/add0/n9730 , \SADR/ADDIDX/add_x_y/add0/n9739 , 
        \SADR/ADDIDX/add_x_y/add0/n9745 , \SADR/ADDIDX/add_x_y/add0/n9737 , 
        \SADR/ADDIDX/add_x_y/add0/n9742 , \SADR/ADDIDX/add_x_y/add0/n9750 , 
        \SADR/ADDIDX/add_x_y/add0/n9736 , \SADR/ADDIDX/add_x_y/add0/n9743 , 
        \SADR/ADDIDX/add_x_y/add0/n9738 , \SADR/ADDIDX/add_x_y/add0/n9751 , 
        \SADR/ADDIDX/add_x_y/add0/n9731 , \SADR/ADDIDX/add_x_y/add0/n9744 , 
        \SADR/ADDIDX/add_x_y/add1/c_last , \SADR/ADDIDX/add_x_y/add1/n9696 , 
        \SADR/ADDIDX/add_x_y/add1/n9706 , \SADR/ADDIDX/add_x_y/add1/n9714 , 
        \SADR/ADDIDX/add_x_y/add1/n9713 , \SADR/ADDIDX/add_x_y/add1/n9688 , 
        \SADR/ADDIDX/add_x_y/add1/n9689 , \SADR/ADDIDX/add_x_y/add1/n9690 , 
        \SADR/ADDIDX/add_x_y/add1/n9691 , \SADR/ADDIDX/add_x_y/add1/n9698 , 
        \SADR/ADDIDX/add_x_y/add1/n9708 , \SADR/ADDIDX/add_x_y/add1/n9699 , 
        \SADR/ADDIDX/add_x_y/add1/n9701 , \SADR/ADDIDX/add_x_y/add1/n9700 , 
        \SADR/ADDIDX/add_x_y/add1/n9709 , \SADR/ADDIDX/add_x_y/add1/n9712 , 
        \SADR/ADDIDX/add_x_y/add1/n9697 , \SADR/ADDIDX/add_x_y/add1/n9707 , 
        \SADR/ADDIDX/add_x_y/add1/n9715 , \SADR/ADDIDX/add_x_y/add1/n9695 , 
        \SADR/ADDIDX/add_x_y/add1/n9705 , \SADR/ADDIDX/add_x_y/add1/n9710 , 
        \SADR/ADDIDX/add_x_y/add1/n9717 , \SADR/ADDIDX/add_x_y/add1/n9719 , 
        \SADR/ADDIDX/add_x_y/add1/n9692 , \SADR/ADDIDX/add_x_y/add1/n9702 , 
        \SADR/ADDIDX/add_x_y/add1/n9693 , \SADR/ADDIDX/add_x_y/add1/n9711 , 
        \SADR/ADDIDX/add_x_y/add1/n9703 , \SADR/ADDIDX/add_x_y/add1/n9694 , 
        \SADR/ADDIDX/add_x_y/add1/n9704 , \SADR/ADDIDX/add_x_y/add1/n9718 , 
        \SADR/ADDIDX/add_x_y/add1/n9716 , \SADR/ADDIDX/add_x_y/add2/c_last , 
        \SADR/ADDIDX/add_x_y/add2/n9668 , \SADR/ADDIDX/add_x_y/add2/n9673 , 
        \SADR/ADDIDX/add_x_y/add2/n9684 , \SADR/ADDIDX/add_x_y/add2/n9661 , 
        \SADR/ADDIDX/add_x_y/add2/n9666 , \SADR/ADDIDX/add_x_y/add2/n9683 , 
        \SADR/ADDIDX/add_x_y/add2/n9656 , \SADR/ADDIDX/add_x_y/add2/n9657 , 
        \SADR/ADDIDX/add_x_y/add2/n9660 , \SADR/ADDIDX/add_x_y/add2/n9667 , 
        \SADR/ADDIDX/add_x_y/add2/n9674 , \SADR/ADDIDX/add_x_y/add2/n9682 , 
        \SADR/ADDIDX/add_x_y/add2/n9669 , \SADR/ADDIDX/add_x_y/add2/n9675 , 
        \SADR/ADDIDX/add_x_y/add2/n9672 , \SADR/ADDIDX/add_x_y/add2/n9685 , 
        \SADR/ADDIDX/add_x_y/add2/n9670 , \SADR/ADDIDX/add_x_y/add2/n9658 , 
        \SADR/ADDIDX/add_x_y/add2/n9659 , \SADR/ADDIDX/add_x_y/add2/n9662 , 
        \SADR/ADDIDX/add_x_y/add2/n9679 , \SADR/ADDIDX/add_x_y/add2/n9687 , 
        \SADR/ADDIDX/add_x_y/add2/n9665 , \SADR/ADDIDX/add_x_y/add2/n9680 , 
        \SADR/ADDIDX/add_x_y/add2/n9677 , \SADR/ADDIDX/add_x_y/add2/n9664 , 
        \SADR/ADDIDX/add_x_y/add2/n9681 , \SADR/ADDIDX/add_x_y/add2/n9671 , 
        \SADR/ADDIDX/add_x_y/add2/n9676 , \SADR/ADDIDX/add_x_y/add2/n9663 , 
        \SADR/ADDIDX/add_x_y/add2/n9678 , \SADR/ADDIDX/add_x_y/add2/n9686 , 
        \SADR/ADDIDX/add_x_y/add3/n9633 , \SADR/ADDIDX/add_x_y/add3/n9654 , 
        \SADR/ADDIDX/add_x_y/add3/n9628 , \SADR/ADDIDX/add_x_y/add3/n9641 , 
        \SADR/ADDIDX/add_x_y/add3/n9646 , \SADR/ADDIDX/add_x_y/add3/n9624 , 
        \SADR/ADDIDX/add_x_y/add3/n9625 , \SADR/ADDIDX/add_x_y/add3/n9626 , 
        \SADR/ADDIDX/add_x_y/add3/n9634 , \SADR/ADDIDX/add_x_y/add3/n9648 , 
        \SADR/ADDIDX/add_x_y/add3/n9627 , \SADR/ADDIDX/add_x_y/add3/n9635 , 
        \SADR/ADDIDX/add_x_y/add3/n9653 , \SADR/ADDIDX/add_x_y/add3/n9640 , 
        \SADR/ADDIDX/add_x_y/add3/n9652 , \SADR/ADDIDX/add_x_y/add3/n9649 , 
        \SADR/ADDIDX/add_x_y/add3/n9647 , \SADR/ADDIDX/add_x_y/add3/n9655 , 
        \SADR/ADDIDX/add_x_y/add3/n9629 , \SADR/ADDIDX/add_x_y/add3/n9630 , 
        \SADR/ADDIDX/add_x_y/add3/n9632 , \SADR/ADDIDX/add_x_y/add3/n9639 , 
        \SADR/ADDIDX/add_x_y/add3/n9637 , \SADR/ADDIDX/add_x_y/add3/n9642 , 
        \SADR/ADDIDX/add_x_y/add3/n9645 , \SADR/ADDIDX/add_x_y/add3/n9636 , 
        \SADR/ADDIDX/add_x_y/add3/n9650 , \SADR/ADDIDX/add_x_y/add3/n9643 , 
        \SADR/ADDIDX/add_x_y/add3/n9651 , \SADR/ADDIDX/add_x_y/add3/n9631 , 
        \SADR/ADDIDX/add_x_y/add3/n9638 , \SADR/ADDIDX/add_x_y/add3/n9644 , 
        \SADR/ADDIDX/add_w_x_z/add0/c_last , 
        \SADR/ADDIDX/add_w_x_z/add0/n9593 , \SADR/ADDIDX/add_w_x_z/add0/n9606 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9621 , \SADR/ADDIDX/add_w_x_z/add0/n9614 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9594 , \SADR/ADDIDX/add_w_x_z/add0/n9591 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9592 , 
        \SADR/ADDIDX/add_w_x_z/add0/gp_out , 
        \SADR/ADDIDX/add_w_x_z/add0/n9595 , \SADR/ADDIDX/add_w_x_z/add0/n9601 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9608 , \SADR/ADDIDX/add_w_x_z/add0/n9613 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9612 , \SADR/ADDIDX/add_w_x_z/add0/n9600 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9609 , \SADR/ADDIDX/add_w_x_z/add0/n9607 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9620 , \SADR/ADDIDX/add_w_x_z/add0/n9596 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9597 , \SADR/ADDIDX/add_w_x_z/add0/n9615 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9599 , \SADR/ADDIDX/add_w_x_z/add0/n9605 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9622 , \SADR/ADDIDX/add_w_x_z/add0/n9617 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9602 , \SADR/ADDIDX/add_w_x_z/add0/n9610 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9611 , \SADR/ADDIDX/add_w_x_z/add0/n9619 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9598 , \SADR/ADDIDX/add_w_x_z/add0/n9603 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9618 , \SADR/ADDIDX/add_w_x_z/add0/n9604 , 
        \SADR/ADDIDX/add_w_x_z/add0/n9616 , 
        \SADR/ADDIDX/add_w_x_z/add1/c_last , 
        \SADR/ADDIDX/add_w_x_z/add1/n9564 , \SADR/ADDIDX/add_w_x_z/add1/n9581 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9588 , \SADR/ADDIDX/add_w_x_z/add1/n9571 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9576 , \SADR/ADDIDX/add_w_x_z/add1/n9559 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9562 , \SADR/ADDIDX/add_w_x_z/add1/n9563 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9578 , \SADR/ADDIDX/add_w_x_z/add1/n9586 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9570 , \SADR/ADDIDX/add_w_x_z/add1/n9579 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9587 , \SADR/ADDIDX/add_w_x_z/add1/n9560 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9565 , \SADR/ADDIDX/add_w_x_z/add1/n9580 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9577 , \SADR/ADDIDX/add_w_x_z/add1/n9589 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9567 , \SADR/ADDIDX/add_w_x_z/add1/n9569 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9572 , \SADR/ADDIDX/add_w_x_z/add1/n9575 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9582 , \SADR/ADDIDX/add_w_x_z/add1/n9590 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9585 , \SADR/ADDIDX/add_w_x_z/add1/n9561 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9568 , \SADR/ADDIDX/add_w_x_z/add1/n9573 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9566 , \SADR/ADDIDX/add_w_x_z/add1/n9583 , 
        \SADR/ADDIDX/add_w_x_z/add1/n9584 , \SADR/ADDIDX/add_w_x_z/add1/n9574 , 
        \SADR/ADDIDX/add_w_x_z/add2/c_last , 
        \SADR/ADDIDX/add_w_x_z/add2/n9536 , \SADR/ADDIDX/add_w_x_z/add2/n9543 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9558 , \SADR/ADDIDX/add_w_x_z/add2/n9551 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9556 , \SADR/ADDIDX/add_w_x_z/add2/n9527 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9530 , \SADR/ADDIDX/add_w_x_z/add2/n9531 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9538 , \SADR/ADDIDX/add_w_x_z/add2/n9539 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9544 , \SADR/ADDIDX/add_w_x_z/add2/n9545 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9557 , \SADR/ADDIDX/add_w_x_z/add2/n9537 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9542 , \SADR/ADDIDX/add_w_x_z/add2/n9550 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9535 , \SADR/ADDIDX/add_w_x_z/add2/n9540 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9549 , \SADR/ADDIDX/add_w_x_z/add2/n9528 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9529 , \SADR/ADDIDX/add_w_x_z/add2/n9532 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9552 , \SADR/ADDIDX/add_w_x_z/add2/n9555 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9546 , \SADR/ADDIDX/add_w_x_z/add2/n9547 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9554 , \SADR/ADDIDX/add_w_x_z/add2/n9533 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9534 , \SADR/ADDIDX/add_w_x_z/add2/n9541 , 
        \SADR/ADDIDX/add_w_x_z/add2/n9548 , \SADR/ADDIDX/add_w_x_z/add2/n9553 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9503 , \SADR/ADDIDX/add_w_x_z/add3/n9511 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9524 , \SADR/ADDIDX/add_w_x_z/add3/n9518 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9495 , \SADR/ADDIDX/add_w_x_z/add3/n9504 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9523 , \SADR/ADDIDX/add_w_x_z/add3/n9516 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9522 , \SADR/ADDIDX/add_w_x_z/add3/n9496 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9497 , \SADR/ADDIDX/add_w_x_z/add3/n9505 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9510 , \SADR/ADDIDX/add_w_x_z/add3/n9517 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9499 , \SADR/ADDIDX/add_w_x_z/add3/n9502 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9519 , \SADR/ADDIDX/add_w_x_z/add3/n9525 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9500 , \SADR/ADDIDX/add_w_x_z/add3/n9509 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9512 , \SADR/ADDIDX/add_w_x_z/add3/n9506 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9507 , \SADR/ADDIDX/add_w_x_z/add3/n9515 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9520 , \SADR/ADDIDX/add_w_x_z/add3/n9498 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9508 , \SADR/ADDIDX/add_w_x_z/add3/n9513 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9514 , \SADR/ADDIDX/add_w_x_z/add3/n9521 , 
        \SADR/ADDIDX/add_w_x_z/add3/n9501 , \SADR/ADDIDX/add_w_x_z/add3/n9526 , 
        \SADR/ADDIDX/add_w_y_z/add0/c_last , 
        \SADR/ADDIDX/add_w_y_z/add0/n9464 , \SADR/ADDIDX/add_w_y_z/add0/n9481 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9476 , \SADR/ADDIDX/add_w_y_z/add0/n9493 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9488 , \SADR/ADDIDX/add_w_y_z/add0/n9462 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9463 , \SADR/ADDIDX/add_w_y_z/add0/n9471 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9470 , \SADR/ADDIDX/add_w_y_z/add0/n9478 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9486 , \SADR/ADDIDX/add_w_y_z/add0/n9479 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9487 , 
        \SADR/ADDIDX/add_w_y_z/add0/gp_out , 
        \SADR/ADDIDX/add_w_y_z/add0/n9465 , \SADR/ADDIDX/add_w_y_z/add0/n9480 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9466 , \SADR/ADDIDX/add_w_y_z/add0/n9467 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9477 , \SADR/ADDIDX/add_w_y_z/add0/n9489 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9492 , \SADR/ADDIDX/add_w_y_z/add0/n9482 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9468 , \SADR/ADDIDX/add_w_y_z/add0/n9469 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9475 , \SADR/ADDIDX/add_w_y_z/add0/n9490 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9472 , \SADR/ADDIDX/add_w_y_z/add0/n9473 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9485 , \SADR/ADDIDX/add_w_y_z/add0/n9484 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9474 , \SADR/ADDIDX/add_w_y_z/add0/n9483 , 
        \SADR/ADDIDX/add_w_y_z/add0/n9491 , 
        \SADR/ADDIDX/add_w_y_z/add1/c_last , 
        \SADR/ADDIDX/add_w_y_z/add1/n9436 , \SADR/ADDIDX/add_w_y_z/add1/n9458 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9443 , \SADR/ADDIDX/add_w_y_z/add1/n9451 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9430 , \SADR/ADDIDX/add_w_y_z/add1/n9431 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9438 , \SADR/ADDIDX/add_w_y_z/add1/n9444 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9456 , \SADR/ADDIDX/add_w_y_z/add1/n9439 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9457 , \SADR/ADDIDX/add_w_y_z/add1/n9432 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9437 , \SADR/ADDIDX/add_w_y_z/add1/n9442 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9445 , \SADR/ADDIDX/add_w_y_z/add1/n9459 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9435 , \SADR/ADDIDX/add_w_y_z/add1/n9450 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9440 , \SADR/ADDIDX/add_w_y_z/add1/n9447 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9449 , \SADR/ADDIDX/add_w_y_z/add1/n9452 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9455 , \SADR/ADDIDX/add_w_y_z/add1/n9460 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9433 , \SADR/ADDIDX/add_w_y_z/add1/n9454 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9434 , \SADR/ADDIDX/add_w_y_z/add1/n9441 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9446 , \SADR/ADDIDX/add_w_y_z/add1/n9461 , 
        \SADR/ADDIDX/add_w_y_z/add1/n9448 , \SADR/ADDIDX/add_w_y_z/add1/n9453 , 
        \SADR/ADDIDX/add_w_y_z/add2/c_last , 
        \SADR/ADDIDX/add_w_y_z/add2/n9399 , \SADR/ADDIDX/add_w_y_z/add2/n9411 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9418 , \SADR/ADDIDX/add_w_y_z/add2/n9403 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9424 , \SADR/ADDIDX/add_w_y_z/add2/n9404 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9423 , \SADR/ADDIDX/add_w_y_z/add2/n9398 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9405 , \SADR/ADDIDX/add_w_y_z/add2/n9416 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9410 , \SADR/ADDIDX/add_w_y_z/add2/n9417 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9422 , \SADR/ADDIDX/add_w_y_z/add2/n9402 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9425 , \SADR/ADDIDX/add_w_y_z/add2/n9400 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9419 , \SADR/ADDIDX/add_w_y_z/add2/n9409 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9412 , \SADR/ADDIDX/add_w_y_z/add2/n9401 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9406 , \SADR/ADDIDX/add_w_y_z/add2/n9407 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9420 , \SADR/ADDIDX/add_w_y_z/add2/n9427 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9415 , \SADR/ADDIDX/add_w_y_z/add2/n9429 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9421 , \SADR/ADDIDX/add_w_y_z/add2/n9408 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9414 , \SADR/ADDIDX/add_w_y_z/add2/n9428 , 
        \SADR/ADDIDX/add_w_y_z/add2/n9413 , \SADR/ADDIDX/add_w_y_z/add2/n9426 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9375 , \SADR/ADDIDX/add_w_y_z/add3/n9382 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9390 , \SADR/ADDIDX/add_w_y_z/add3/n9367 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9385 , \SADR/ADDIDX/add_w_y_z/add3/n9366 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9368 , \SADR/ADDIDX/add_w_y_z/add3/n9369 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9372 , \SADR/ADDIDX/add_w_y_z/add3/n9397 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9373 , \SADR/ADDIDX/add_w_y_z/add3/n9384 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9396 , \SADR/ADDIDX/add_w_y_z/add3/n9374 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9391 , \SADR/ADDIDX/add_w_y_z/add3/n9370 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9371 , \SADR/ADDIDX/add_w_y_z/add3/n9383 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9376 , \SADR/ADDIDX/add_w_y_z/add3/n9378 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9381 , \SADR/ADDIDX/add_w_y_z/add3/n9393 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9388 , \SADR/ADDIDX/add_w_y_z/add3/n9386 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9394 , \SADR/ADDIDX/add_w_y_z/add3/n9379 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9387 , \SADR/ADDIDX/add_w_y_z/add3/n9377 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9389 , \SADR/ADDIDX/add_w_y_z/add3/n9395 , 
        \SADR/ADDIDX/add_w_y_z/add3/n9392 , \SADR/ADDIDX/add_w_y_z/add3/n9380 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/c_last , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9335 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9349 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9352 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9340 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9347 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9360 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9333 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9355 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9334 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/gp_out , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9341 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9346 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9348 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9354 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9361 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9353 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9336 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9351 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9358 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9337 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9338 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9343 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9344 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9363 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9364 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9339 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9345 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9356 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9362 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9357 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9342 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9350 , 
        \SADR/ADDIDX/add_w_x_y_z/add0/n9359 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/c_last , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9312 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9327 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9309 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9301 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9306 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9307 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9315 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9329 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9332 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9320 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9314 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9321 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9328 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9302 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9303 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9326 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9308 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9313 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9318 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9324 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9304 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9311 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9316 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9331 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9305 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9317 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9323 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9330 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9322 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9325 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9310 , 
        \SADR/ADDIDX/add_w_x_y_z/add1/n9319 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/c_last , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9275 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9290 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9300 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9282 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9299 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9269 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9272 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9285 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9297 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9270 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9271 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9273 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9284 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9296 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9274 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9291 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9283 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9298 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9276 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9288 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9293 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9278 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9281 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9286 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9279 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9287 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9294 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9295 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9277 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9280 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9289 , 
        \SADR/ADDIDX/add_w_x_y_z/add2/n9292 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9240 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9249 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9252 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9267 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9237 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9238 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9246 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9247 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9260 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9255 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9261 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9248 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9253 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9254 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9268 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9241 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9243 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9266 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9251 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9264 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9244 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9258 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9256 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9263 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9239 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9245 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9262 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9250 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9257 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9259 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9242 , 
        \SADR/ADDIDX/add_w_x_y_z/add3/n9265 , 
        \REGF/pbmemff41/phdec12_2/dec4_1/n7077 , 
        \REGF/pbmemff41/phdec12_2/dec4_1/n7079 , 
        \REGF/pbmemff41/phdec12_2/dec4_1/n7076 , 
        \REGF/pbmemff41/phdec12_2/dec4_1/n7078 , 
        \REGF/pbmemff41/phdec12_2/dec4_1/n7075 , 
        \REGF/pbmemff41/phdec12_2/dec4_3/n7070 , 
        \REGF/pbmemff41/phdec12_2/dec4_3/n7071 , 
        \REGF/pbmemff41/phdec12_2/dec4_3/gg_out , 
        \REGF/pbmemff41/phdec12_2/dec4_3/n7073 , 
        \REGF/pbmemff41/phdec12_2/dec4_3/n7074 , 
        \REGF/pbmemff41/phdec12_2/dec4_3/n7072 , 
        \REGF/pbmemff41/phdec12_2/dec4_2/n7065 , 
        \REGF/pbmemff41/phdec12_2/dec4_2/n7066 , 
        \REGF/pbmemff41/phdec12_2/dec4_2/n7068 , 
        \REGF/pbmemff41/phdec12_2/dec4_2/n7069 , 
        \REGF/pbmemff41/phdec12_2/dec4_2/n7067 , 
        \REGF/pbmemff41/phdec12_1/dec4_1/n7059 , 
        \REGF/pbmemff41/phdec12_1/dec4_1/n7062 , 
        \REGF/pbmemff41/phdec12_1/dec4_1/n7058 , 
        \REGF/pbmemff41/phdec12_1/dec4_1/n7061 , 
        \REGF/pbmemff41/phdec12_1/dec4_1/n7060 , 
        \REGF/pbmemff41/phdec12_1/dec4_3/n7057 , 
        \REGF/pbmemff41/phdec12_1/dec4_3/n7056 , 
        \REGF/pbmemff41/phdec12_1/dec4_3/gg_out , 
        \REGF/pbmemff41/phdec12_1/dec4_3/n7053 , 
        \REGF/pbmemff41/phdec12_1/dec4_3/n7054 , 
        \REGF/pbmemff41/phdec12_1/dec4_3/n7055 , 
        \REGF/pbmemff41/phdec12_1/dec4_2/n7050 , 
        \REGF/pbmemff41/phdec12_1/dec4_2/n7051 , 
        \REGF/pbmemff41/phdec12_1/dec4_2/n7048 , 
        \REGF/pbmemff41/phdec12_1/dec4_2/n7052 , 
        \REGF/pbmemff41/phdec12_1/dec4_2/n7049 , 
        \MAIN/ENGIN/STEP_A/deocgen_1/n3543 , 
        \MAIN/ENGIN/STEP_B/deocgen_1/n3495 , 
        \MAIN/ENGIN/STEP_C/deocgen_1/n3447 , 
        \MAIN/ENGIN/STEP_D/deocgen_1/n3399 , \ALUSHT/ALU/dec32/dec4_7/n1800 , 
        \ALUSHT/ALU/dec32/dec4_7/gg_out , \ALUSHT/ALU/dec32/dec4_7/n1797 , 
        \ALUSHT/ALU/dec32/dec4_7/n1799 , \ALUSHT/ALU/dec32/dec4_7/n1798 , 
        \ALUSHT/ALU/dec32/dec4_7/n1796 , \ALUSHT/ALU/dec32/dec4_0/n1793 , 
        \ALUSHT/ALU/dec32/dec4_0/n1794 , \ALUSHT/ALU/dec32/dec4_0/n1792 , 
        \ALUSHT/ALU/dec32/dec4_0/n1795 , \ALUSHT/ALU/dec32/dec4_0/n1791 , 
        \ALUSHT/ALU/dec32/dec4_1/n1786 , \ALUSHT/ALU/dec32/dec4_1/n1788 , 
        \ALUSHT/ALU/dec32/dec4_1/n1789 , \ALUSHT/ALU/dec32/dec4_1/n1787 , 
        \ALUSHT/ALU/dec32/dec4_1/n1790 , \ALUSHT/ALU/dec32/dec4_2/n1781 , 
        \ALUSHT/ALU/dec32/dec4_2/n1785 , \ALUSHT/ALU/dec32/dec4_2/n1782 , 
        \ALUSHT/ALU/dec32/dec4_2/n1783 , \ALUSHT/ALU/dec32/dec4_2/n1784 , 
        \ALUSHT/ALU/dec32/dec4_3/n1778 , \ALUSHT/ALU/dec32/dec4_3/n1776 , 
        \ALUSHT/ALU/dec32/dec4_3/n1777 , \ALUSHT/ALU/dec32/dec4_3/n1779 , 
        \ALUSHT/ALU/dec32/dec4_3/n1780 , \ALUSHT/ALU/dec32/dec4_4/n1771 , 
        \ALUSHT/ALU/dec32/dec4_4/n1772 , \ALUSHT/ALU/dec32/dec4_4/n1775 , 
        \ALUSHT/ALU/dec32/dec4_4/n1774 , \ALUSHT/ALU/dec32/dec4_4/n1773 , 
        \ALUSHT/ALU/dec32/dec4_6/n1770 , \ALUSHT/ALU/dec32/dec4_6/n1767 , 
        \ALUSHT/ALU/dec32/dec4_6/n1769 , \ALUSHT/ALU/dec32/dec4_6/n1766 , 
        \ALUSHT/ALU/dec32/dec4_6/n1768 , \ALUSHT/ALU/dec32/dec4_5/n1763 , 
        \ALUSHT/ALU/dec32/dec4_5/n1636 , \ALUSHT/ALU/dec32/dec4_5/n1764 , 
        \ALUSHT/ALU/dec32/dec4_5/n1637 , \ALUSHT/ALU/dec32/dec4_5/n1765 , 
        \ALUSHT/ALU/add32/add0/c_last , \ALUSHT/ALU/add32/add0/n1359 , 
        \ALUSHT/ALU/add32/add0/n1365 , \ALUSHT/ALU/add32/add0/n1377 , 
        \ALUSHT/ALU/add32/add0/n1380 , \ALUSHT/ALU/add32/add0/n1357 , 
        \ALUSHT/ALU/add32/add0/n1358 , \ALUSHT/ALU/add32/add0/n1362 , 
        \ALUSHT/ALU/add32/add0/n1370 , \ALUSHT/ALU/add32/add0/n1387 , 
        \ALUSHT/ALU/add32/add0/n1363 , \ALUSHT/ALU/add32/add0/n1371 , 
        \ALUSHT/ALU/add32/add0/n1379 , \ALUSHT/ALU/add32/add0/n1378 , 
        \ALUSHT/ALU/add32/add0/n1364 , \ALUSHT/ALU/add32/add0/n1381 , 
        \ALUSHT/ALU/add32/add0/n1386 , \ALUSHT/ALU/add32/add0/n1388 , 
        \ALUSHT/ALU/add32/add0/n1360 , \ALUSHT/ALU/add32/add0/n1361 , 
        \ALUSHT/ALU/add32/add0/n1376 , \ALUSHT/ALU/add32/add0/n1366 , 
        \ALUSHT/ALU/add32/add0/n1368 , \ALUSHT/ALU/add32/add0/n1374 , 
        \ALUSHT/ALU/add32/add0/n1383 , \ALUSHT/ALU/add32/add0/n1373 , 
        \ALUSHT/ALU/add32/add0/n1384 , \ALUSHT/ALU/add32/add0/n1369 , 
        \ALUSHT/ALU/add32/add0/n1372 , \ALUSHT/ALU/add32/add0/n1367 , 
        \ALUSHT/ALU/add32/add0/n1382 , \ALUSHT/ALU/add32/add0/n1385 , 
        \ALUSHT/ALU/add32/add0/n1375 , \ALUSHT/ALU/add32/add1/c_last , 
        \ALUSHT/ALU/add32/add1/n1337 , \ALUSHT/ALU/add32/add1/n1342 , 
        \ALUSHT/ALU/add32/add1/n1350 , \ALUSHT/ALU/add32/add1/n1325 , 
        \ALUSHT/ALU/add32/add1/n1326 , \ALUSHT/ALU/add32/add1/n1330 , 
        \ALUSHT/ALU/add32/add1/n1339 , \ALUSHT/ALU/add32/add1/n1345 , 
        \ALUSHT/ALU/add32/add1/n1331 , \ALUSHT/ALU/add32/add1/n1338 , 
        \ALUSHT/ALU/add32/add1/n1356 , \ALUSHT/ALU/add32/add1/n1336 , 
        \ALUSHT/ALU/add32/add1/n1343 , \ALUSHT/ALU/add32/add1/n1344 , 
        \ALUSHT/ALU/add32/add1/n1351 , \ALUSHT/ALU/add32/add1/n1334 , 
        \ALUSHT/ALU/add32/add1/n1341 , \ALUSHT/ALU/add32/add1/n1348 , 
        \ALUSHT/ALU/add32/add1/n1353 , \ALUSHT/ALU/add32/add1/n1327 , 
        \ALUSHT/ALU/add32/add1/n1328 , \ALUSHT/ALU/add32/add1/n1354 , 
        \ALUSHT/ALU/add32/add1/n1329 , \ALUSHT/ALU/add32/add1/n1332 , 
        \ALUSHT/ALU/add32/add1/n1333 , \ALUSHT/ALU/add32/add1/n1346 , 
        \ALUSHT/ALU/add32/add1/n1355 , \ALUSHT/ALU/add32/add1/n1347 , 
        \ALUSHT/ALU/add32/add1/n1335 , \ALUSHT/ALU/add32/add1/n1340 , 
        \ALUSHT/ALU/add32/add1/n1349 , \ALUSHT/ALU/add32/add1/n1352 , 
        \ALUSHT/ALU/add32/add2/c_last , \ALUSHT/ALU/add32/add2/n1310 , 
        \ALUSHT/ALU/add32/add2/n1319 , \ALUSHT/ALU/add32/add2/n1295 , 
        \ALUSHT/ALU/add32/add2/n1302 , \ALUSHT/ALU/add32/add2/n1305 , 
        \ALUSHT/ALU/add32/add2/n1322 , \ALUSHT/ALU/add32/add2/n1293 , 
        \ALUSHT/ALU/add32/add2/n1294 , \ALUSHT/ALU/add32/add2/n1317 , 
        \ALUSHT/ALU/add32/add2/n1323 , \ALUSHT/ALU/add32/add2/n1303 , 
        \ALUSHT/ALU/add32/add2/n1304 , \ALUSHT/ALU/add32/add2/n1311 , 
        \ALUSHT/ALU/add32/add2/n1316 , \ALUSHT/ALU/add32/add2/n1296 , 
        \ALUSHT/ALU/add32/add2/n1298 , \ALUSHT/ALU/add32/add2/n1324 , 
        \ALUSHT/ALU/add32/add2/n1318 , \ALUSHT/ALU/add32/add2/n1313 , 
        \ALUSHT/ALU/add32/add2/n1301 , \ALUSHT/ALU/add32/add2/n1308 , 
        \ALUSHT/ALU/add32/add2/n1297 , \ALUSHT/ALU/add32/add2/n1306 , 
        \ALUSHT/ALU/add32/add2/n1307 , \ALUSHT/ALU/add32/add2/n1314 , 
        \ALUSHT/ALU/add32/add2/n1321 , \ALUSHT/ALU/add32/add2/n1299 , 
        \ALUSHT/ALU/add32/add2/n1309 , \ALUSHT/ALU/add32/add2/n1315 , 
        \ALUSHT/ALU/add32/add2/n1320 , \ALUSHT/ALU/add32/add2/n1300 , 
        \ALUSHT/ALU/add32/add2/n1312 , \ALUSHT/ALU/add32/add5/n1280 , 
        \ALUSHT/ALU/add32/add5/n1289 , \ALUSHT/ALU/add32/add5/n1277 , 
        \ALUSHT/ALU/add32/add5/n1292 , \ALUSHT/ALU/add32/add5/n1273 , 
        \ALUSHT/ALU/add32/add5/n1274 , \ALUSHT/ALU/add32/add5/n1278 , 
        \ALUSHT/ALU/add32/add5/n1279 , \ALUSHT/ALU/add32/add5/n1287 , 
        \ALUSHT/ALU/add32/add5/n1286 , \ALUSHT/ALU/add32/add5/n1281 , 
        \ALUSHT/ALU/add32/add5/n1276 , \ALUSHT/ALU/add32/add5/n1288 , 
        \ALUSHT/ALU/add32/add5/n1283 , \ALUSHT/ALU/add32/add5/n1291 , 
        \ALUSHT/ALU/add32/add5/n1275 , \ALUSHT/ALU/add32/add5/n1282 , 
        \ALUSHT/ALU/add32/add5/n1284 , \ALUSHT/ALU/add32/add5/n1285 , 
        \ALUSHT/ALU/add32/add5/n1290 , \ALUSHT/ALU/add32/add3/c_last , 
        \ALUSHT/ALU/add32/add3/n1242 , \ALUSHT/ALU/add32/add3/n1259 , 
        \ALUSHT/ALU/add32/add3/n1265 , \ALUSHT/ALU/add32/add3/n1250 , 
        \ALUSHT/ALU/add32/add3/n1270 , \ALUSHT/ALU/add32/add3/n1241 , 
        \ALUSHT/ALU/add32/add3/n1243 , \ALUSHT/ALU/add32/add3/n1244 , 
        \ALUSHT/ALU/add32/add3/n1245 , \ALUSHT/ALU/add32/add3/n1257 , 
        \ALUSHT/ALU/add32/add3/n1262 , \ALUSHT/ALU/add32/add3/n1256 , 
        \ALUSHT/ALU/add32/add3/n1271 , \ALUSHT/ALU/add32/add3/n1263 , 
        \ALUSHT/ALU/add32/add3/n1258 , \ALUSHT/ALU/add32/add3/n1264 , 
        \ALUSHT/ALU/add32/add3/n1251 , \ALUSHT/ALU/add32/add3/n1266 , 
        \ALUSHT/ALU/add32/add3/n1246 , \ALUSHT/ALU/add32/add3/n1248 , 
        \ALUSHT/ALU/add32/add3/n1253 , \ALUSHT/ALU/add32/add3/n1254 , 
        \ALUSHT/ALU/add32/add3/n1268 , \ALUSHT/ALU/add32/add3/n1247 , 
        \ALUSHT/ALU/add32/add3/n1255 , \ALUSHT/ALU/add32/add3/n1261 , 
        \ALUSHT/ALU/add32/add3/n1269 , \ALUSHT/ALU/add32/add3/n1272 , 
        \ALUSHT/ALU/add32/add3/n1249 , \ALUSHT/ALU/add32/add3/n1252 , 
        \ALUSHT/ALU/add32/add3/n1260 , \ALUSHT/ALU/add32/add3/n1267 , 
        \ALUSHT/ALU/add32/add4/c_last , \ALUSHT/ALU/add32/add4/n1225 , 
        \ALUSHT/ALU/add32/add4/n1237 , \ALUSHT/ALU/add32/add4/n1239 , 
        \ALUSHT/ALU/add32/add4/n1221 , \ALUSHT/ALU/add32/add4/n1222 , 
        \ALUSHT/ALU/add32/add4/n1223 , \ALUSHT/ALU/add32/add4/n1230 , 
        \ALUSHT/ALU/add32/add4/n1231 , \ALUSHT/ALU/add32/add4/n1238 , 
        \ALUSHT/ALU/add32/add4/n1236 , \ALUSHT/ALU/add32/add4/n1224 , 
        \ALUSHT/ALU/add32/add4/n1226 , \ALUSHT/ALU/add32/add4/n1234 , 
        \ALUSHT/ALU/add32/add4/n1227 , \ALUSHT/ALU/add32/add4/n1228 , 
        \ALUSHT/ALU/add32/add4/n1233 , \ALUSHT/ALU/add32/add4/n1229 , 
        \ALUSHT/ALU/add32/add4/n1232 , \ALUSHT/ALU/add32/add4/n1235 , 
        \ALUSHT/ALU/add32/add4/n1240 , \ALUSHT/ALU/cmp32/cmp4_7/n1197 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1202 , \ALUSHT/ALU/cmp32/cmp4_7/n1210 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1199 , \ALUSHT/ALU/cmp32/cmp4_7/n1205 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1194 , \ALUSHT/ALU/cmp32/cmp4_7/n1196 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1198 , \ALUSHT/ALU/cmp32/cmp4_7/n1204 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1203 , \ALUSHT/ALU/cmp32/cmp4_7/n1208 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1201 , \ALUSHT/ALU/cmp32/cmp4_7/n1206 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1207 , \ALUSHT/ALU/cmp32/cmp4_7/n1195 , 
        \ALUSHT/ALU/cmp32/cmp4_7/n1209 , \ALUSHT/ALU/cmp32/cmp4_7/n1200 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1182 , \ALUSHT/ALU/cmp32/cmp4_6/n1185 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1177 , \ALUSHT/ALU/cmp32/cmp4_6/n1178 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1183 , \ALUSHT/ALU/cmp32/cmp4_6/n1190 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1191 , \ALUSHT/ALU/cmp32/cmp4_6/n1184 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1180 , \ALUSHT/ALU/cmp32/cmp4_6/n1181 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1186 , \ALUSHT/ALU/cmp32/cmp4_6/n1188 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1193 , \ALUSHT/ALU/cmp32/cmp4_6/n1192 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1189 , \ALUSHT/ALU/cmp32/cmp4_6/n1179 , 
        \ALUSHT/ALU/cmp32/cmp4_6/n1187 , \ALUSHT/ALU/cmp32/cmp4_1/n1169 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1172 , \ALUSHT/ALU/cmp32/cmp4_1/n1160 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1171 , \ALUSHT/ALU/cmp32/cmp4_1/n1175 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1167 , \ALUSHT/ALU/cmp32/cmp4_1/n1161 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1166 , \ALUSHT/ALU/cmp32/cmp4_1/n1168 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1174 , \ALUSHT/ALU/cmp32/cmp4_1/n1173 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1176 , \ALUSHT/ALU/cmp32/cmp4_1/n1163 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1164 , \ALUSHT/ALU/cmp32/cmp4_1/n1165 , 
        \ALUSHT/ALU/cmp32/cmp4_1/n1170 , \ALUSHT/ALU/cmp32/cmp4_1/n1162 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1150 , \ALUSHT/ALU/cmp32/cmp4_0/n1155 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1147 , \ALUSHT/ALU/cmp32/cmp4_0/n1156 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1152 , \ALUSHT/ALU/cmp32/cmp4_0/n1149 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1154 , \ALUSHT/ALU/cmp32/cmp4_0/n1153 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1148 , \ALUSHT/ALU/cmp32/cmp4_0/n1146 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1158 , \ALUSHT/ALU/cmp32/cmp4_0/n1143 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1144 , \ALUSHT/ALU/cmp32/cmp4_0/n1159 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1151 , \ALUSHT/ALU/cmp32/cmp4_0/n1157 , 
        \ALUSHT/ALU/cmp32/cmp4_0/n1145 , \ALUSHT/ALU/cmp32/cmp4_5/n1132 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1129 , \ALUSHT/ALU/cmp32/cmp4_5/n1127 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1135 , \ALUSHT/ALU/cmp32/cmp4_5/n1140 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1126 , \ALUSHT/ALU/cmp32/cmp4_5/n1134 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1141 , \ALUSHT/ALU/cmp32/cmp4_5/n1128 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1131 , \ALUSHT/ALU/cmp32/cmp4_5/n1133 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1138 , \ALUSHT/ALU/cmp32/cmp4_5/n1136 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1137 , \ALUSHT/ALU/cmp32/cmp4_5/n1142 , 
        \ALUSHT/ALU/cmp32/cmp4_5/n1130 , \ALUSHT/ALU/cmp32/cmp4_5/n1139 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1115 , \ALUSHT/ALU/cmp32/cmp4_4/n1120 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1109 , \ALUSHT/ALU/cmp32/cmp4_4/n1112 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1110 , \ALUSHT/ALU/cmp32/cmp4_4/n1111 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1113 , \ALUSHT/ALU/cmp32/cmp4_4/n1114 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1121 , \ALUSHT/ALU/cmp32/cmp4_4/n1116 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1123 , \ALUSHT/ALU/cmp32/cmp4_4/n1118 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1124 , \ALUSHT/ALU/cmp32/cmp4_4/n1119 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1122 , \ALUSHT/ALU/cmp32/cmp4_4/n1125 , 
        \ALUSHT/ALU/cmp32/cmp4_4/n1117 , \ALUSHT/ALU/cmp32/cmp4_3/n1099 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1097 , \ALUSHT/ALU/cmp32/cmp4_3/n1107 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1105 , \ALUSHT/ALU/cmp32/cmp4_3/n1106 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1100 , \ALUSHT/ALU/cmp32/cmp4_3/n1096 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1098 , \ALUSHT/ALU/cmp32/cmp4_3/n1101 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1108 , \ALUSHT/ALU/cmp32/cmp4_3/n1093 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1094 , \ALUSHT/ALU/cmp32/cmp4_3/n1103 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1104 , \ALUSHT/ALU/cmp32/cmp4_3/n1092 , 
        \ALUSHT/ALU/cmp32/cmp4_3/n1102 , \ALUSHT/ALU/cmp32/cmp4_3/n1095 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1085 , \ALUSHT/ALU/cmp32/cmp4_2/n1082 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1090 , \ALUSHT/ALU/cmp32/cmp4_2/n1078 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1083 , \ALUSHT/ALU/cmp32/cmp4_2/n1084 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1091 , \ALUSHT/ALU/cmp32/cmp4_2/n1086 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1080 , \ALUSHT/ALU/cmp32/cmp4_2/n1081 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1088 , \ALUSHT/ALU/cmp32/cmp4_2/n1089 , 
        \ALUSHT/ALU/cmp32/cmp4_2/n1079 , \ALUSHT/ALU/cmp32/cmp4_2/n1087 , 
        \ALUSHT/ALU/inc32/inc4_0/n1075 , \ALUSHT/ALU/inc32/inc4_0/n1076 , 
        \ALUSHT/ALU/inc32/inc4_0/n1077 , \ALUSHT/ALU/inc32/inc4_1/n1072 , 
        \ALUSHT/ALU/inc32/inc4_1/n1073 , \ALUSHT/ALU/inc32/inc4_1/n1074 , 
        \ALUSHT/ALU/inc32/inc4_6/n1069 , \ALUSHT/ALU/inc32/inc4_6/n1071 , 
        \ALUSHT/ALU/inc32/inc4_6/n1070 , \ALUSHT/ALU/inc32/inc4_7/gp_out , 
        \ALUSHT/ALU/inc32/inc4_7/n1066 , \ALUSHT/ALU/inc32/inc4_7/n1067 , 
        \ALUSHT/ALU/inc32/inc4_7/n1068 , \ALUSHT/ALU/inc32/inc4_2/n1063 , 
        \ALUSHT/ALU/inc32/inc4_2/n1064 , \ALUSHT/ALU/inc32/inc4_2/n1065 , 
        \ALUSHT/ALU/inc32/inc4_3/n1060 , \ALUSHT/ALU/inc32/inc4_3/n1061 , 
        \ALUSHT/ALU/inc32/inc4_3/n1062 , \ALUSHT/ALU/inc32/inc4_4/n1058 , 
        \ALUSHT/ALU/inc32/inc4_4/n1059 , \ALUSHT/ALU/inc32/inc4_4/n1057 , 
        \ALUSHT/ALU/inc32/inc4_5/n1055 , \ALUSHT/ALU/inc32/inc4_5/n1052 , 
        \ALUSHT/ALU/inc32/inc4_5/n1053 , \ALUSHT/ALU/inc32/inc4_5/n1054 , 
        \ALUSHT/ALU/inc32/inc4_5/n1056 ;
    assign PDH[63] = SWIT_wire;
    assign PDH[62] = SWIT_wire;
    assign PDH[61] = SWIT_wire;
    assign PDH[60] = SWIT_wire;
    assign SWIT_wire = SWIT;
    snl_invx1 U4 ( .ZN(n10737), .A(phrstihb) );
    snl_invx1 U5 ( .ZN(n10732), .A(n10737) );
    snl_invx1 U6 ( .ZN(n10731), .A(n10737) );
    snl_bufx1 \REGF/U376  ( .Z(\REGF/n8052 ), .A(n10732) );
    snl_oai222x2 \REGF/U388  ( .ZN(\REGF/RI_SRA12M[24] ), .A(\REGF/n8065 ), 
        .B(\REGF/n8051 ), .C(\REGF/n8227 ), .D(\REGF/n8158 ), .E(\REGF/n8228 ), 
        .F(\REGF/n8157 ) );
    snl_ao022x1 \REGF/U409  ( .Z(\REGF/RI_PCOH[24] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[24]), .C(\stream4[56] ), .D(\REGF/n8053 ) );
    snl_oai012x1 \LBUS/U563  ( .ZN(LTC0), .A(word32odtrh), .B(ph_locken_h), 
        .C(\LBUS/ilt[2] ) );
    snl_oai222x0 \REGF/U440  ( .ZN(\REGF/RI_EACC[25] ), .A(\REGF/n8073 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8074 ), .E(\REGF/n8075 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U482  ( .ZN(\REGF/RI_DPR[11] ), .A(\REGF/n8185 ), .B(
        \REGF/n8160 ), .C(\REGF/n8186 ), .D(\REGF/n8162 ), .E(\REGF/n8117 ), 
        .F(\REGF/n8151 ) );
    snl_oai222x0 \REGF/U599  ( .ZN(\REGF/RI_ACC[2] ), .A(\REGF/n8142 ), .B(
        \REGF/n8215 ), .C(\REGF/n8143 ), .D(\REGF/n8216 ), .E(\REGF/n8144 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U739  ( .ZN(\REGF/n8085 ), .A(\pgldi[21] ) );
    snl_invx05 \CODEIF/U265  ( .ZN(\CODEIF/n3879 ), .A(PDLIN[4]) );
    snl_xnor2x0 \CONS/U214  ( .ZN(\CONS/n701 ), .A(\pk_pc_h[9] ), .B(
        \pk_pcs1_h[9] ) );
    snl_nor03x0 \BLU/U403  ( .ZN(\BLU/n1574 ), .A(all0bsel), .B(accbsel), .C(
        srcbsel) );
    snl_and02x1 \REG_2/U145  ( .Z(\ph_cpudout[15] ), .A(\ph_segset_h[15] ), 
        .B(seg_cnfg_h) );
    snl_invx05 \BLU/U382  ( .ZN(\BLU/n1506 ), .A(\pgld16[2] ) );
    snl_oai122x0 \ADOSEL/U19  ( .ZN(\pgmuxout[8] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4113 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4114 ), .E(
        \ADOSEL/n4115 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[0]  ( .Q(\CODEIF/pfctr[0] ), .D(
        \CODEIF/pfctr415[0] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_muxi21x1 \LDIS/U193  ( .ZN(\LDIS/ldexch[17] ), .A(\LDIS/n3150 ), .B(
        \LDIS/n3149 ), .S(\LDIS/n3165 ) );
    snl_aoi123x0 \LBUS/U653  ( .ZN(\LBUS/n1429 ), .A(\LBUS/n1600 ), .B(LDK), 
        .C(\LBUS/n1424 ), .D(\LBUS/n1605 ), .E(\LBUS/n1417 ), .F(ph_d53lth) );
    snl_nor02x1 \PDOSEL/U128  ( .ZN(\PDOSEL/n183 ), .A(\pk_pdo_h[15] ), .B(
        \ph_cpudout[15] ) );
    snl_nand03x0 \LBUS/U674  ( .ZN(\LBUS/n1442 ), .A(\LBUS/ilt[0] ), .B(
        \LBUS/n1456 ), .C(\LBUS/n1460 ) );
    snl_xor2x0 \CONS/U86  ( .Z(\CONS/n604 ), .A(\pk_idcz_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_and08x1 \CONS/U124  ( .Z(\CONS/n558 ), .A(\CONS/n649 ), .B(\CONS/n650 
        ), .C(\CONS/n651 ), .D(\CONS/n652 ), .E(\CONS/n653 ), .F(\CONS/n654 ), 
        .G(\CONS/n655 ), .H(\CONS/n648 ) );
    snl_nor02x1 \CODEIF/U242  ( .ZN(\CODEIF/n3928 ), .A(\CODEIF/n3926 ), .B(
        \CODEIF/wprotect1 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[13]  ( .Q(\CODEIF/pfctr[13] ), .D(
        \CODEIF/pfctr415[13] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_xor2x0 \CONS/U103  ( .Z(\CONS/n621 ), .A(\pk_idcx_h[19] ), .B(
        \pk_indx_h[19] ) );
    snl_invx05 \REG_2/U162  ( .ZN(\REG_2/n517 ), .A(ph_initldh) );
    snl_and02x1 \ALUIS/U27  ( .Z(\ALUIS/n3655 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3665 ) );
    snl_and02x1 \LDIS/U228  ( .Z(\LDIS/n3134 ), .A(ph_word32_h), .B(
        \pgsadrh[1] ) );
    snl_xnor2x0 \CONS/U233  ( .ZN(\CONS/n720 ), .A(\pk_idcy_h[5] ), .B(
        \pk_indy_h[5] ) );
    snl_invx05 \BLU/U424  ( .ZN(\BLU/n1528 ), .A(\BLU/n1480 ) );
    snl_oai022x1 \BLU/U309  ( .ZN(\pkbludgh[7] ), .A(\BLU/n1464 ), .B(
        \BLU/n1489 ), .C(\BLU/n1490 ), .D(\BLU/n1491 ) );
    snl_ao022x1 \REGF/U512  ( .Z(\REGF/RI_PCOL[13] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[13]), .C(\stream4[13] ), .D(\REGF/n8209 ) );
    snl_ao2222x1 \REGF/U535  ( .Z(\REGF/RI_SRDA[22] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[22]), .C(\pgldi[22] ), .D(\REGF/n8210 ), .E(\stream3[22] ), .F(
        \REGF/n8211 ), .G(\pkdptout[22] ), .H(\REGF/n8212 ) );
    snl_oai022x1 \REGF/U605  ( .ZN(\REGF/RI_SPR[24] ), .A(\REGF/n8157 ), .B(
        \REGF/n8218 ), .C(\REGF/n8219 ), .D(\REGF/n8158 ) );
    snl_oai222x0 \REGF/U622  ( .ZN(\REGF/RI_SPR[7] ), .A(\REGF/n8193 ), .B(
        \REGF/n8220 ), .C(\REGF/n8194 ), .D(\REGF/n8221 ), .E(\REGF/n8129 ), 
        .F(\REGF/n8218 ) );
    snl_oai022x1 \MAIN/U171  ( .ZN(\MAIN/n3624 ), .A(\MAIN/c_exec_stage ), .B(
        ph_dec_dh), .C(\MAIN/a_exec_stage ), .D(ph_dec_bh) );
    snl_xor2x0 \LDCHK/U64  ( .Z(\LDCHK/n3294 ), .A(\pgld32[7] ), .B(
        \pgld32[2] ) );
    snl_ao022x1 \LDIS/U118  ( .Z(\pgldi[10] ), .A(ph_word32_h), .B(
        \pgld32[10] ), .C(\pgld16[10] ), .D(ph_word16_h) );
    snl_nand02x1 \ADOSEL/U92  ( .ZN(\ADOSEL/n4151 ), .A(\pgbluext[28] ), .B(
        \ADOSEL/n4156 ) );
    snl_invx05 \MAIN/U156  ( .ZN(\MAIN/n3623 ), .A(\MAIN/n3626 ) );
    snl_xnor2x0 \CONS/U188  ( .ZN(\CONS/n669 ), .A(\pgsdprlh[21] ), .B(
        \CONS/SACO[17] ) );
    snl_ao022x1 \BLUOS/U19  ( .Z(\pgbluext[31] ), .A(\pkbludgh[15] ), .B(
        ph_bit_h), .C(\pkdptout[15] ), .D(ph_word16_h) );
    snl_invx05 \REGF/U795  ( .ZN(\REGF/n8068 ), .A(\pkdptout[27] ) );
    snl_xor2x0 \CODEIF/U359  ( .Z(\CODEIF/n3935 ), .A(CDIN[31]), .B(
        \CODEIF/n3949 ) );
    snl_nor03x0 \LDCHK/U43  ( .ZN(\LDCHK/n3240 ), .A(\pgld32[29] ), .B(
        \pgld32[30] ), .C(\LDCHK/n3255 ) );
    snl_nand02x1 \ALUIS/U169  ( .ZN(\ALUIS/n3673 ), .A(\pk_ada_h[15] ), .B(
        po_arsel_h) );
    snl_invx05 \REGF/U770  ( .ZN(\REGF/n8172 ), .A(\pgsdprlh[18] ) );
    snl_nand02x1 \ADOSEL/U108  ( .ZN(\ADOSEL/n4130 ), .A(\pgbluext[29] ), .B(
        \ADOSEL/n4156 ) );
    snl_ao222x1 \CODEIF/U197  ( .Z(\CODEIF/n3844 ), .A(PA[6]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[3] ), .E(cif_byte), .F(PDLIN[3])
         );
    snl_invx05 \LDIS/U151  ( .ZN(\LDIS/n3120 ), .A(\pgld32[20] ) );
    snl_oai012x1 \PDOSEL/U35  ( .ZN(PDH[51]), .A(\PDOSEL/n105 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_xor2x0 \CODEIF/U337  ( .Z(\CODEIF/n4020 ), .A(CDOUT[14]), .B(CDOUT[4])
         );
    snl_or02x1 \MAIN/U138  ( .Z(\MAIN/sprw_inhibith ), .A(\MAIN/sprw_tap2 ), 
        .B(\MAIN/sprw_tap1 ) );
    snl_mux21x1 \ALUSHT/U22  ( .Z(\pkdptout[29] ), .A(\ALUSHT/pkshtout[29] ), 
        .B(\ALUSHT/pkaluout[29] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U63  ( .Z(\CONS/n580 ), .A(\CONS/SACO[4] ), .B(
        \pgsdprlh[8] ) );
    snl_nor02x1 \SAEXE/U106  ( .ZN(ph_srcadr1_h), .A(\SAEXE/n417 ), .B(
        \SAEXE/n413 ) );
    snl_oai112x0 \LBUS/U691  ( .ZN(\LBUS/n1606 ), .A(\LBUS/temp[3] ), .B(
        \LBUS/n1452 ), .C(\LBUS/ilt[0] ), .D(\LBUS/ilt[1] ) );
    snl_invx05 \BLU/U340  ( .ZN(\BLU/n1555 ), .A(\poalufnc[2] ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[13]  ( .Q(CA[13]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3854 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_aoi022x1 \ALUIS/U107  ( .ZN(\ALUIS/n3742 ), .A(\stream4[26] ), .B(
        immbsel), .C(\pk_adb_h[26] ), .D(po_brsel_h) );
    snl_invx05 \CODEIF/U280  ( .ZN(\CODEIF/n3908 ), .A(\CODEIF/pfctr[14] ) );
    snl_xor2x0 \CODEIF/U310  ( .Z(\CODEIF/n3953 ), .A(\CODEIF/n3980 ), .B(
        \CODEIF/n3981 ) );
    snl_nand02x1 \ALUIS/U49  ( .ZN(\pgaluinb[1] ), .A(\ALUIS/n3692 ), .B(
        \ALUIS/n3693 ) );
    snl_invx05 \LDCHK/U122  ( .ZN(\LDCHK/n3308 ), .A(\pgld32[26] ) );
    snl_aoi012x1 \ALUIS/U120  ( .ZN(\ALUIS/n3693 ), .A(\pgldi[1] ), .B(srcbsel
        ), .C(allfbsel) );
    snl_xnor2x0 \LDCHK/U105  ( .ZN(\LDCHK/n3282 ), .A(\pgmuxout[18] ), .B(
        \pgmuxout[17] ) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[6]  ( .Q(\REG_2/RETCNT[6] ), .D(
        \REG_2/ph_retcnt_h[6] ), .EN(\REG_2/n517 ), .RN(\REG_2/n436 ), .SD(
        \REG_2/ncnt3[0] ), .SE(ph_d76lth), .CP(SCLK) );
    snl_nor04x0 \BLU/U367  ( .ZN(\BLU/n1572 ), .A(\BLU/n1550 ), .B(\BLU/n1544 
        ), .C(\BLU/n1549 ), .D(\BLU/n1531 ) );
    snl_ffqx1 \LDCHK/pchkenh_reg  ( .Q(\LDCHK/pchkenh ), .D(LPDIN), .CP(SCLK)
         );
    snl_muxi21x1 \LDIS/U176  ( .ZN(\LDIS/ldexcl[11] ), .A(\LDIS/n3159 ), .B(
        \LDIS/n3160 ), .S(\LDIS/n3134 ) );
    snl_and02x1 \LBUS/U586  ( .Z(ph_lbe3_h), .A(\LBUS/EXTSEL ), .B(phsaerrh)
         );
    snl_nand13x1 \CONS/U44  ( .ZN(\CONS/n550 ), .A(word32odtrh), .B(
        \pk_saco_lh[4] ), .C(ph_lwdsrc_h) );
    snl_aoi012x1 \SAEXE/U121  ( .ZN(\SAEXE/n417 ), .A(\SAEXE/n430 ), .B(
        \SAEXE/n422 ), .C(\SAEXE/rf_srcadr1_h ) );
    snl_invx05 \ADOSEL/U77  ( .ZN(\ADOSEL/n4092 ), .A(\pkdptout[17] ) );
    snl_ffqrnx1 \CODEIF/pgpaendp_reg  ( .Q(pgpaendp), .D(\CODEIF/frpend_in ), 
        .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nand02x1 \PDOSEL/U161  ( .ZN(\PDOSEL/n126 ), .A(CDIN[11]), .B(
        \PDOSEL/n119 ) );
    snl_oai022x1 \REGF/U467  ( .ZN(\REGF/RI_DPR[26] ), .A(\REGF/n8062 ), .B(
        \REGF/n8151 ), .C(\REGF/n8152 ), .D(\REGF/n8154 ) );
    snl_muxi21x1 \REGF/U832  ( .ZN(\REGF/n8231 ), .A(\REGF/n8239 ), .B(
        \REGF/n8234 ), .S(\REGF/RO_ACC[17] ) );
    snl_and02x1 \REGF/U567  ( .Z(\REGF/RO_LPSAS2156[9] ), .A(ph_sastlth), .B(
        ph_byrtendh) );
    snl_and02x1 \REGF/U657  ( .Z(pkaccovf), .A(\REGF/n8231 ), .B(po_raccen_h)
         );
    snl_invx05 \REGF/U757  ( .ZN(\REGF/n8198 ), .A(\pgsdprlh[5] ) );
    snl_nor04x0 \REGF/U815  ( .ZN(\REGF/n8234 ), .A(\REGF/n8235 ), .B(
        \REGF/n8236 ), .C(\REGF/n8237 ), .D(\REGF/n8238 ) );
    snl_aoi022x1 \LDCHK/U81  ( .ZN(\LDCHK/n3307 ), .A(\LDCHK/n3308 ), .B(
        \LDCHK/n3239 ), .C(\pgld32[26] ), .D(\pgld32[27] ) );
    snl_and02x1 \REGF/U829  ( .Z(\REGF/n8227 ), .A(\REGF/n8229 ), .B(
        \REGF/n8230 ) );
    snl_invx05 \ADOSEL/U50  ( .ZN(\ADOSEL/n4110 ), .A(\pkdptout[23] ) );
    snl_invx05 \PDOSEL/U99  ( .ZN(\PDOSEL/n101 ), .A(CDIN[47]) );
    snl_ao222x1 \CODEIF/U210  ( .Z(\CODEIF/n3857 ), .A(PA[19]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[16] ), .E(cif_byte), .F(PDLIN[16]
        ) );
    snl_xnor2x0 \CODEIF/U380  ( .ZN(\CODEIF/n3975 ), .A(CDIN[35]), .B(CDIN[34]
        ) );
    snl_invx1 \ALUIS/U9  ( .ZN(\pgaluina[10] ), .A(\ALUIS/n3641 ) );
    snl_ao022x1 \LDIS/U98  ( .Z(\pgldi[0] ), .A(ph_word32_h), .B(\pgld32[0] ), 
        .C(\pgld16[0] ), .D(ph_word16_h) );
    snl_nand02x1 \PDOSEL/U146  ( .ZN(\PDOSEL/n148 ), .A(CDIN[24]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \PDOSEL/U82  ( .ZN(\PDOSEL/n81 ), .A(CDIN[37]) );
    snl_sffqenrnx1 \LDCHK/pglpinff_reg[0]  ( .Q(\LDCHK/pglpinff[0] ), .D(1'b0), 
        .EN(1'b1), .RN(n10733), .SD(\LDCHK/lpex[0] ), .SE(ph_lpdilth), .CP(
        SCLK) );
    snl_nand03x0 \CONS/U151  ( .ZN(\CONS/n722 ), .A(\CONS/n723 ), .B(
        \CONS/n724 ), .C(\CONS/n725 ) );
    snl_nor02x1 \LBUS/U626  ( .ZN(\LBUS/n1596 ), .A(\LBUS/n1595 ), .B(
        ph_errtendh) );
    snl_ao022x1 \REG_2/U130  ( .Z(\ph_cpudout[0] ), .A(\ph_segset_h[0] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[0] ), .D(ret_cont_h) );
    snl_xnor2x0 \CODEIF/U401  ( .ZN(\CODEIF/n3995 ), .A(CDOUT[58]), .B(CDOUT
        [59]) );
    snl_xnor2x0 \CONS/U261  ( .ZN(\CONS/n743 ), .A(\pk_idcw_h[11] ), .B(
        \pk_indw_h[11] ) );
    snl_oai122x0 \CODEIF/U237  ( .ZN(\CODEIF/pfctr415[16] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3914 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3915 ), .E(
        \CODEIF/n3916 ) );
    snl_xnor2x0 \CONS/U246  ( .ZN(\CONS/n731 ), .A(\pk_idcx_h[5] ), .B(
        \pk_indx_h[5] ) );
    snl_aoi112x0 \LBUS/U601  ( .ZN(\LBUS/n1408 ), .A(ph_lbslock_h), .B(
        \LBUS/n1404 ), .C(\LBUS/n1454 ), .D(\LBUS/n1436 ) );
    snl_xnor2x0 \CONS/U176  ( .ZN(\CONS/n655 ), .A(\pgsdprlh[5] ), .B(
        \pk_saco_lh[5] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[7]  ( .Q(\ph_segset_h[7] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[7]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_nand02x3 \REGF/U393  ( .ZN(\REGF/n8216 ), .A(ph_rgfile_h), .B(
        \REGF/n8217 ) );
    snl_ao022x1 \REGF/U412  ( .Z(\REGF/RI_PCOH[21] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[21]), .C(\stream4[53] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U435  ( .ZN(\REGF/RI_EACC[30] ), .A(\REGF/n8060 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8061 ), .E(\REGF/n8062 ), 
        .F(\REGF/n8059 ) );
    snl_ao022x1 \REGF/U499  ( .Z(\REGF/RI_PCOL[26] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[26]), .C(\stream4[26] ), .D(\REGF/n8209 ) );
    snl_ao2222x1 \REGF/U540  ( .Z(\REGF/RI_SRDA[17] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[17]), .C(\pgldi[17] ), .D(\REGF/n8210 ), .E(\stream3[17] ), .F(
        \REGF/n8211 ), .G(\pkdptout[17] ), .H(\REGF/n8212 ) );
    snl_nand02x1 \ALUIS/U52  ( .ZN(\pgaluinb[4] ), .A(\ALUIS/n3698 ), .B(
        \ALUIS/n3699 ) );
    snl_oai022x1 \REGF/U639  ( .ZN(\REGF/RI_TBAI[18] ), .A(\REGF/n8225 ), .B(
        \REGF/n8084 ), .C(\REGF/n8226 ), .D(\REGF/n8163 ) );
    snl_invx05 \REGF/U670  ( .ZN(\REGF/n8191 ), .A(\pgregadrh[8] ) );
    snl_nand02x1 \ALUIS/U75  ( .ZN(\pgaluinb[27] ), .A(\ALUIS/n3744 ), .B(
        \ALUIS/n3745 ) );
    snl_and08x1 \LDCHK/U36  ( .A(\LDCHK/n3238 ), .B(\LDCHK/n3239 ), .C(
        \LDCHK/n3240 ), .D(\LDCHK/n3241 ), .E(\LDCHK/n3230 ), .F(\LDCHK/n3242 
        ), .G(\LDCHK/n3243 ), .H(\LDCHK/n3244 ) );
    snl_mux21x1 \ALUSHT/U39  ( .Z(\pkdptout[13] ), .A(\ALUSHT/pkshtout[13] ), 
        .B(\ALUSHT/pkaluout[13] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U78  ( .Z(\CONS/n596 ), .A(\pk_pcs1_h[15] ), .B(
        \pk_pc_h[15] ) );
    snl_nand02x1 \CODEIF/U342  ( .ZN(\CODEIF/n3886 ), .A(\CODEIF/pgctrinc[6] ), 
        .B(\CODEIF/n3945 ) );
    snl_nand02x1 \MAIN/U123  ( .ZN(\MAIN/*cell*4603/U14/CONTROL1 ), .A(
        \MAIN/n3613 ), .B(\MAIN/n3615 ) );
    snl_nand02x1 \ALUIS/U172  ( .ZN(\ALUIS/n3670 ), .A(\pk_ada_h[12] ), .B(
        po_arsel_h) );
    snl_nand02x1 \ADOSEL/U89  ( .ZN(\ADOSEL/n4153 ), .A(\pgbluext[30] ), .B(
        \ADOSEL/n4156 ) );
    snl_xor2x0 \LDCHK/U58  ( .Z(\LDCHK/n3258 ), .A(\LDCHK/n3282 ), .B(
        \LDCHK/n3283 ) );
    snl_invx05 \LDIS/U214  ( .ZN(\LDIS/n3133 ), .A(LIN[25]) );
    snl_nor02x1 \BLU/U335  ( .ZN(\BLU/n1478 ), .A(\BLU/n1532 ), .B(\BLU/n1550 
        ) );
    snl_ao022x1 \LDIS/U124  ( .Z(\pgldi[13] ), .A(ph_word32_h), .B(
        \pgld32[13] ), .C(\pgld16[13] ), .D(ph_word16_h) );
    snl_ffandx1 \LBUS/lnsa_end_reg  ( .Q(\LBUS/lnsa_end ), .A(\LBUS/temp[3] ), 
        .B(\LBUS/*cell*3982/U158/Z_0 ), .CP(SCLK) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[9]  ( .Q(\CODEIF/pfctr[9] ), .D(
        \CODEIF/pfctr415[9] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_xnor2x0 \CONS/U193  ( .ZN(\CONS/n681 ), .A(\pk_pc_h[8] ), .B(
        \pk_pcs2_h[8] ) );
    snl_oai012x1 \PDOSEL/U40  ( .ZN(PDH[56]), .A(\PDOSEL/n110 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_ao022x1 \BLUOS/U25  ( .Z(\pgbluext[6] ), .A(\pkbludgh[6] ), .B(
        ph_bit_h), .C(\pkdptout[6] ), .D(ph_word16_h) );
    snl_and08x1 \CONS/U31  ( .Z(ph_izco_h), .A(\CONS/n528 ), .B(\CONS/n529 ), 
        .C(\CONS/n530 ), .D(\CONS/n531 ), .E(\CONS/n532 ), .F(\CONS/n533 ), 
        .G(\CONS/n534 ), .H(\CONS/n535 ) );
    snl_ao022x1 \LDIS/U103  ( .Z(\pgld16[2] ), .A(ph_selldl), .B(\pgld32[2] ), 
        .C(ph_selldh), .D(\pgld32[18] ) );
    snl_or02x1 \CMPX/U12  ( .Z(ph_lbussth), .A(phrelbsth), .B(lbus_start) );
    snl_oai112x0 \PDOSEL/U67  ( .ZN(PDLOUT[6]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n82 ), .C(\PDOSEL/n156 ), .D(\PDOSEL/n157 ) );
    snl_ao022x1 \REGF/U509  ( .Z(\REGF/RI_PCOL[16] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[16]), .C(\stream4[16] ), .D(\REGF/n8209 ) );
    snl_invx05 \CODEIF/U259  ( .ZN(\CODEIF/n3888 ), .A(PDLIN[7]) );
    snl_xor2x0 \CODEIF/U365  ( .Z(\CODEIF/n4026 ), .A(\CODEIF/n4027 ), .B(
        \CODEIF/n4013 ) );
    snl_oai022x1 \BLU/U312  ( .ZN(\pkbludgh[4] ), .A(\BLU/n1464 ), .B(
        \BLU/n1498 ), .C(\BLU/n1499 ), .D(\BLU/n1500 ) );
    snl_aoi012x1 \ALUIS/U90  ( .ZN(\ALUIS/n3699 ), .A(\pgldi[4] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_nand02x1 \ALUIS/U155  ( .ZN(\ALUIS/n3686 ), .A(\pk_ada_h[28] ), .B(
        po_arsel_h) );
    snl_xnor2x0 \CONS/U228  ( .ZN(\CONS/n529 ), .A(\pk_idcz_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_invx05 \REGF/U695  ( .ZN(\REGF/n8093 ), .A(PDLIN[19]) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[6]  ( .Q(CA[6]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3847 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_xor2x0 \CONS/U118  ( .Z(\CONS/n636 ), .A(\pk_idcw_h[22] ), .B(
        \pk_indw_h[22] ) );
    snl_nor02x1 \PDOSEL/U114  ( .ZN(\PDOSEL/n145 ), .A(\pk_pdo_h[2] ), .B(
        \ph_cpudout[2] ) );
    snl_invx05 \REGF/U705  ( .ZN(\REGF/n8108 ), .A(PDLIN[14]) );
    snl_invx05 \REGF/U722  ( .ZN(\REGF/n8141 ), .A(PDLIN[3]) );
    snl_oai122x0 \ADOSEL/U25  ( .ZN(\pgmuxout[14] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4131 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4132 ), .E(
        \ADOSEL/n4133 ) );
    snl_nor02x1 \PDOSEL/U133  ( .ZN(\PDOSEL/n116 ), .A(\ph_cpudout[10] ), .B(
        \pk_pdo_h[10] ) );
    snl_muxi21x1 \LDIS/U188  ( .ZN(\LDIS/ldexch[22] ), .A(\LDIS/n3140 ), .B(
        \LDIS/n3139 ), .S(\LDIS/n3165 ) );
    snl_aoi022x1 \LBUS/U648  ( .ZN(\LBUS/n1591 ), .A(\LBUS/n1452 ), .B(
        \LBUS/n1456 ), .C(\LBUS/ilt[4] ), .D(\LBUS/ilt[1] ) );
    snl_nand02x1 \BLU/U399  ( .ZN(\BLU/n1480 ), .A(\BLU/n1562 ), .B(
        \BLU/n1561 ) );
    snl_invx05 \BLU/U418  ( .ZN(\BLU/n1543 ), .A(\BLU/n1504 ) );
    snl_ao022x1 \REGF/U427  ( .Z(\REGF/RI_PCOH[6] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[6]), .C(\stream4[38] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U582  ( .ZN(\REGF/RI_ACC[19] ), .A(\REGF/n8091 ), .B(
        \REGF/n8215 ), .C(\REGF/n8092 ), .D(\REGF/n8216 ), .E(\REGF/n8093 ), 
        .F(\REGF/n8217 ) );
    snl_aoi012x1 \ALUIS/U82  ( .ZN(\ALUIS/n3707 ), .A(\pgldi[8] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_and34x0 \LBUS/U578  ( .Z(ph_sprlth), .A(\LBUS/n1438 ), .B(\LBUS/n1439 
        ), .C(\LBUS/n1406 ), .D(po_sprlth) );
    snl_invx05 \REGF/U687  ( .ZN(\REGF/n8081 ), .A(PDLIN[23]) );
    snl_invx05 \REGF/U717  ( .ZN(\REGF/n8127 ), .A(\pgldi[7] ) );
    snl_invx1 \ADOSEL/U10  ( .ZN(\ADOSEL/n4156 ), .A(ph_word32_h) );
    snl_nor04x0 \PDOSEL/U106  ( .ZN(\PDOSEL/n225 ), .A(BE[0]), .B(BE[3]), .C(
        BE[2]), .D(BE[1]) );
    snl_oai122x0 \ADOSEL/U37  ( .ZN(\pgmuxout[26] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4120 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4119 ), .E(
        \ADOSEL/n4149 ) );
    snl_oai2222x0 \REGF/U364  ( .ZN(\REGF/RI_SRA12M[6] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8132 ), .C(\REGF/n8130 ), .D(\REGF/n8051 ), .E(\REGF/n8195 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8196 ) );
    snl_oai2222x0 \REGF/U381  ( .ZN(\REGF/RI_SRA12M[16] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8102 ), .C(\REGF/n8100 ), .D(\REGF/n8051 ), .E(\REGF/n8175 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8176 ) );
    snl_invx1 \REGF/U400  ( .ZN(\REGF/n8218 ), .A(\ph_pdis_h[3] ) );
    snl_oai222x0 \REGF/U590  ( .ZN(\REGF/RI_ACC[11] ), .A(\REGF/n8115 ), .B(
        \REGF/n8215 ), .C(\REGF/n8116 ), .D(\REGF/n8216 ), .E(\REGF/n8117 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U730  ( .ZN(\REGF/n8069 ), .A(PDLIN[27]) );
    snl_nor02x1 \PDOSEL/U121  ( .ZN(\PDOSEL/n159 ), .A(\pk_pdo_h[21] ), .B(
        \ph_cpudout[21] ) );
    snl_oai022x1 \REGF/U645  ( .ZN(\REGF/RI_TBAI[12] ), .A(\REGF/n8225 ), .B(
        \REGF/n8102 ), .C(\REGF/n8226 ), .D(\REGF/n8175 ) );
    snl_nand02x1 \CODEIF/U350  ( .ZN(\CODEIF/n3916 ), .A(\CODEIF/pgctrinc[16] 
        ), .B(\CODEIF/n3945 ) );
    snl_invx05 \LDIS/U206  ( .ZN(\LDIS/n3142 ), .A(LIN[21]) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[2]  ( .Q(\REG_2/RETCNT[2] ), .D(
        \REG_2/ph_retcnt_h[2] ), .EN(\REG_2/n517 ), .RN(\REG_2/n436 ), .SD(
        \REG_2/ncnt1[2] ), .SE(ph_d20lth), .CP(SCLK) );
    snl_nor04x0 \BLU/U327  ( .ZN(\BLU/n1499 ), .A(\BLU/n1535 ), .B(\BLU/n1537 
        ), .C(\BLU/n1538 ), .D(\BLU/n1534 ) );
    snl_nand02x1 \ALUIS/U160  ( .ZN(\ALUIS/n3681 ), .A(\pk_ada_h[23] ), .B(
        po_arsel_h) );
    snl_xor2x0 \CODEIF/U377  ( .Z(\CODEIF/n3931 ), .A(\CODEIF/n3971 ), .B(
        \CODEIF/n4031 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[17]  ( .Q(CA[17]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3858 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_ao022x1 \LDIS/U111  ( .Z(\pgld16[6] ), .A(ph_selldl), .B(\pgld32[6] ), 
        .C(ph_selldh), .D(\pgld32[22] ) );
    snl_oai012x1 \LDIS/U136  ( .ZN(\pgldi[22] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3122 ), .C(\LDIS/n3115 ) );
    snl_ao022x1 \CMPX/U27  ( .Z(ph_bit_h), .A(ph_bitsrch), .B(ph_saexe_sth), 
        .C(srctype0), .D(\CMPX/n1047 ) );
    snl_xnor2x0 \CONS/U181  ( .ZN(\CONS/n657 ), .A(\pgsdprlh[17] ), .B(
        \pk_saco_lh[17] ) );
    snl_oai112x0 \PDOSEL/U52  ( .ZN(PDLOUT[3]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n79 ), .C(\PDOSEL/n128 ), .D(\PDOSEL/n129 ) );
    snl_ffqsnx1 \LBUS/cmd_oe_h_reg  ( .Q(LCMDCNT), .D(\LBUS/n_2434 ), .SN(
        n10734), .CP(SCLK) );
    snl_oai112x0 \PDOSEL/U75  ( .ZN(PDLOUT[15]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n101 ), .C(\PDOSEL/n182 ), .D(\PDOSEL/n183 ) );
    snl_invx05 \LDIS/U221  ( .ZN(\LDIS/n3155 ), .A(LIN[13]) );
    snl_nand02x1 \ALUIS/U147  ( .ZN(\ALUIS/n3664 ), .A(\pk_ada_h[6] ), .B(
        po_arsel_h) );
    snl_muxi21x2 \BLU/U300  ( .ZN(\BLU/n1464 ), .A(\BLU/n1553 ), .B(pk_rgbit_h
        ), .S(ph_dregsl_h) );
    snl_invx05 \SAEXE/U128  ( .ZN(\SAEXE/n429 ), .A(\pk_psae_h[7] ) );
    snl_sffqsnx1 \LBUS/ph_lpdoeh_reg  ( .Q(LPDCNT), .D(\LBUS/n_2439 ), .SN(
        n10734), .SD(\LBUS/n_2434 ), .SE(ph_lbwrh), .CP(SCLK) );
    snl_ao2222x1 \REGF/U552  ( .Z(\REGF/RI_SRDA[5] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[5]), .C(\pgldi[5] ), .D(\REGF/n8210 ), .E(\stream3[5] ), .F(
        \REGF/n8211 ), .G(\pkdptout[5] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U575  ( .ZN(\REGF/RI_ACC[26] ), .A(\REGF/n8070 ), .B(
        \REGF/n8215 ), .C(\REGF/n8071 ), .D(\REGF/n8216 ), .E(\REGF/n8072 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \CODEIF/U289  ( .ZN(\CODEIF/n3897 ), .A(PDLIN[10]) );
    snl_xor2x0 \CODEIF/U319  ( .Z(\CODEIF/n3994 ), .A(\CODEIF/n3995 ), .B(
        \CODEIF/n3996 ) );
    snl_nand02x1 \ALUIS/U40  ( .ZN(\pgaluina[24] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3682 ) );
    snl_aoi022x1 \ALUIS/U129  ( .ZN(\ALUIS/n3722 ), .A(\stream4[16] ), .B(
        immbsel), .C(\pk_adb_h[16] ), .D(po_brsel_h) );
    snl_or02x1 \UPIF/U12  ( .Z(\UPIF/iready ), .A(polcore_end), .B(pgpaendp)
         );
    snl_invx05 \REGF/U662  ( .ZN(\REGF/n8183 ), .A(\pgregadrh[12] ) );
    snl_nand02x1 \ADOSEL/U101  ( .ZN(\ADOSEL/n4094 ), .A(\pgbluext[1] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U67  ( .ZN(\pgaluinb[19] ), .A(\ALUIS/n3728 ), .B(
        \ALUIS/n3729 ) );
    snl_invx05 \BLU/U349  ( .ZN(\BLU/n1564 ), .A(\pgbitnoh[0] ) );
    snl_invx05 \ADOSEL/U59  ( .ZN(\ADOSEL/n4099 ), .A(\pkdptout[3] ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[17]  ( .Q(\CODEIF/pfctr[17] ), .D(
        \CODEIF/pfctr415[17] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_or03x1 \MAIN/U131  ( .Z(\MAIN/EXCEP_EXT ), .A(\MAIN/excep_valid ), .B(
        \MAIN/EXCEP_2H ), .C(\MAIN/EXCEP_1H ) );
    snl_invx05 \LDIS/U158  ( .ZN(\LDIS/n3128 ), .A(\pgld32[28] ) );
    snl_nor03x0 \CONS/U143  ( .ZN(\CONS/n702 ), .A(\CONS/n603 ), .B(
        \CONS/n601 ), .C(\CONS/n602 ) );
    snl_invx05 \PDOSEL/U90  ( .ZN(\PDOSEL/n109 ), .A(CDIN[55]) );
    snl_ao222x1 \CODEIF/U202  ( .Z(\CODEIF/n3849 ), .A(PA[11]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[8] ), .E(cif_byte), .F(PDLIN[8])
         );
    snl_ffqrnx1 \CODEIF/pfctr_reg[4]  ( .Q(\CODEIF/pfctr[4] ), .D(
        \CODEIF/pfctr415[4] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_invx05 \LDCHK/U88  ( .ZN(\LDCHK/n3272 ), .A(LPIN[3]) );
    snl_nor03x0 \LBUS/U634  ( .ZN(\LBUS/n1600 ), .A(\LBUS/ph_lbusylth ), .B(
        LBER), .C(LDS) );
    snl_xor2x0 \CODEIF/U392  ( .Z(\CODEIF/n3956 ), .A(\CODEIF/n4034 ), .B(
        \CODEIF/n4033 ) );
    snl_xnor2x0 \CONS/U273  ( .ZN(\CONS/n339 ), .A(\pk_idcw_h[2] ), .B(
        \pk_indw_h[2] ) );
    snl_xnor2x0 \CODEIF/U413  ( .ZN(\CODEIF/n4009 ), .A(CDOUT[23]), .B(CDOUT
        [28]) );
    snl_sffqenrnx1 \LBUS/word32odtrh_reg  ( .Q(word32odtrh), .D(1'b0), .EN(
        1'b1), .RN(n10734), .SD(\LBUS/*cell*3982/U71/CONTROL1 ), .SE(
        \LBUS/*cell*3982/U148/CONTROL1 ), .CP(SCLK) );
    snl_oai222x0 \REGF/U449  ( .ZN(\REGF/RI_EACC[16] ), .A(\REGF/n8100 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8101 ), .E(\REGF/n8102 ), 
        .F(\REGF/n8059 ) );
    snl_oai122x0 \CODEIF/U225  ( .ZN(\CODEIF/pfctr415[4] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3878 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3879 ), .E(
        \CODEIF/n3880 ) );
    snl_xnor2x0 \CONS/U254  ( .ZN(\CONS/n737 ), .A(\pk_idcx_h[23] ), .B(
        \pk_indx_h[23] ) );
    snl_nand02x1 \BLU/U443  ( .ZN(\BLU/n1580 ), .A(ebaccsel), .B(\BLU/n1553 )
         );
    snl_oai222x0 \REGF/U452  ( .ZN(\REGF/RI_EACC[13] ), .A(\REGF/n8109 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8110 ), .E(\REGF/n8111 ), 
        .F(\REGF/n8059 ) );
    snl_invx05 \REGF/U762  ( .ZN(\REGF/n8203 ), .A(\pgregadrh[2] ) );
    snl_invx05 \REGF/U779  ( .ZN(\REGF/n8208 ), .A(\pgsdprlh[0] ) );
    snl_nand03x0 \LBUS/U613  ( .ZN(\LBUS/n1463 ), .A(\LBUS/ilt[0] ), .B(LDS), 
        .C(\LBUS/ilt[1] ) );
    snl_sffqenrnx1 \LBUS/ph_exstgb_h_reg  ( .Q(ph_exstgb_h), .D(1'b0), .EN(
        1'b1), .RN(n10734), .SD(\LBUS/*cell*3982/U119/CONTROL1 ), .SE(
        \LBUS/*cell*3982/U201/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CONS/U164  ( .ZN(\CONS/n541 ), .A(\CONS/n559 ) );
    snl_or04x1 \REGF/U820  ( .Z(\REGF/n8242 ), .A(\REGF/RO_ACC[27] ), .B(
        \REGF/RO_ACC[20] ), .C(\REGF/RO_ACC[22] ), .D(\REGF/RO_ACC[23] ) );
    snl_invx05 \ADOSEL/U65  ( .ZN(\ADOSEL/n4132 ), .A(\pkdptout[14] ) );
    snl_invx05 \LBUS/U608  ( .ZN(\LBUS/n1456 ), .A(\LBUS/ilt[1] ) );
    snl_oai222x0 \REGF/U475  ( .ZN(\REGF/RI_DPR[18] ), .A(\REGF/n8171 ), .B(
        \REGF/n8160 ), .C(\REGF/n8172 ), .D(\REGF/n8162 ), .E(\REGF/n8096 ), 
        .F(\REGF/n8151 ) );
    snl_invx05 \REGF/U807  ( .ZN(\REGF/n8101 ), .A(\pkdptout[16] ) );
    snl_mux21x1 \SHTCD/U13  ( .Z(\phshtd[4] ), .A(\pgld16[4] ), .B(
        \stream4[4] ), .S(immbsel) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[2]  ( .Q(CA[2]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3843 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_invx05 \REGF/U745  ( .ZN(\REGF/n8100 ), .A(\pgldi[16] ) );
    snl_invx05 \CODEIF/U219  ( .ZN(\CODEIF/n3860 ), .A(n10731) );
    snl_xnor2x0 \CONS/U268  ( .ZN(\CONS/n747 ), .A(\pk_idcw_h[4] ), .B(
        \pk_indw_h[4] ) );
    snl_and02x1 \REG_2/U139  ( .Z(\ph_cpudout[9] ), .A(seg_cnfg_h), .B(
        \ph_segset_h[9] ) );
    snl_xnor2x0 \CODEIF/U389  ( .ZN(\CODEIF/n3954 ), .A(CDIN[22]), .B(CDIN[23]
        ) );
    snl_xnor2x0 \CODEIF/U408  ( .ZN(\CODEIF/n4003 ), .A(CDOUT[43]), .B(CDOUT
        [44]) );
    snl_invx05 \LDCHK/U93  ( .ZN(\LDCHK/n3238 ), .A(\pgld32[0] ) );
    snl_invx2 U7 ( .ZN(n10734), .A(n10737) );
    snl_invx1 U8 ( .ZN(n10733), .A(n10737) );
    snl_ffqx1 \RSTGN/WRST_1H_reg  ( .Q(\RSTGN/WRST_1H ), .D(WRST), .CP(SCLK)
         );
    snl_ffqx1 \RSTGN/CRST_2H_reg  ( .Q(\RSTGN/CRST_2H ), .D(\RSTGN/CRST_1H ), 
        .CP(SCLK) );
    snl_oai2222x0 \REGF/U358  ( .ZN(\REGF/RI_SRA12M[17] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8099 ), .C(\REGF/n8097 ), .D(\REGF/n8051 ), .E(\REGF/n8173 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8174 ) );
    snl_ao2222x1 \REGF/U549  ( .Z(\REGF/RI_SRDA[8] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[8]), .C(\pgldi[8] ), .D(\REGF/n8210 ), .E(\stream3[8] ), .F(
        \REGF/n8211 ), .G(\pkdptout[8] ), .H(\REGF/n8212 ) );
    snl_invx05 \REGF/U679  ( .ZN(\REGF/n8062 ), .A(PDLIN[30]) );
    snl_oai122x0 \ADOSEL/U42  ( .ZN(\pgmuxout[31] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4135 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4134 ), .E(
        \ADOSEL/n4154 ) );
    snl_nand02x1 \PDOSEL/U154  ( .ZN(\PDOSEL/n160 ), .A(CDIN[18]), .B(
        \PDOSEL/n119 ) );
    snl_oai012x1 \LDIS/U143  ( .ZN(\pgldi[29] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3129 ), .C(\LDIS/n3115 ) );
    snl_nor03x0 \CONS/U158  ( .ZN(\CONS/n738 ), .A(\CONS/n630 ), .B(
        \CONS/n628 ), .C(\CONS/n629 ) );
    snl_oai012x1 \PDOSEL/U27  ( .ZN(PDH[43]), .A(\PDOSEL/n97 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_mux21x1 \ALUSHT/U30  ( .Z(\pkdptout[21] ), .A(\ALUSHT/pkshtout[21] ), 
        .B(\ALUSHT/pkaluout[21] ), .S(\ALUSHT/n3112 ) );
    snl_nor02x1 \LBUS/U683  ( .ZN(\LBUS/n1395 ), .A(word32odtrh), .B(
        ph_lbussth) );
    snl_xor2x0 \CONS/U71  ( .Z(\CONS/n589 ), .A(\pk_pcs2_h[13] ), .B(
        \pk_pc_h[13] ) );
    snl_oai022x1 \SAEXE/U114  ( .ZN(phatchkh), .A(\SAEXE/n423 ), .B(
        \SAEXE/n413 ), .C(\SAEXE/n415 ), .D(\SAEXE/n425 ) );
    snl_xor2x0 \CODEIF/U325  ( .Z(\CODEIF/n4004 ), .A(CDOUT[34]), .B(CDOUT[37]
        ) );
    snl_aoi022x1 \ALUIS/U115  ( .ZN(\ALUIS/n3734 ), .A(\stream4[22] ), .B(
        immbsel), .C(\pk_adb_h[22] ), .D(po_brsel_h) );
    snl_nor02x1 \BLU/U352  ( .ZN(\BLU/n1567 ), .A(\BLU/n1566 ), .B(\BLU/n1559 
        ) );
    snl_oai222x0 \REGF/U455  ( .ZN(\REGF/RI_EACC[10] ), .A(\REGF/n8118 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8119 ), .E(\REGF/n8120 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U472  ( .ZN(\REGF/RI_DPR[21] ), .A(\REGF/n8165 ), .B(
        \REGF/n8160 ), .C(\REGF/n8166 ), .D(\REGF/n8162 ), .E(\REGF/n8087 ), 
        .F(\REGF/n8151 ) );
    snl_oai222x0 \REGF/U490  ( .ZN(\REGF/RI_DPR[3] ), .A(\REGF/n8201 ), .B(
        \REGF/n8160 ), .C(\REGF/n8202 ), .D(\REGF/n8162 ), .E(\REGF/n8141 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U500  ( .Z(\REGF/RI_PCOL[25] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[25]), .C(\stream4[25] ), .D(\REGF/n8209 ) );
    snl_xor2x0 \CODEIF/U292  ( .Z(\CODEIF/n3949 ), .A(\CODEIF/n3950 ), .B(
        \CODEIF/n3951 ) );
    snl_xor2x0 \CODEIF/U302  ( .Z(\CODEIF/n3969 ), .A(CDIN[49]), .B(CDIN[48])
         );
    snl_nand02x1 \BLU/U375  ( .ZN(\BLU/n1495 ), .A(\BLU/n1570 ), .B(
        \BLU/n1569 ) );
    snl_nand02x1 \ALUIS/U35  ( .ZN(\pgaluina[19] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3677 ) );
    snl_aoi012x1 \ALUIS/U132  ( .ZN(\ALUIS/n3719 ), .A(\pgldi[14] ), .B(
        srcbsel), .C(allfbsel) );
    snl_aoi022x1 \LDCHK/U117  ( .ZN(\LDCHK/n3310 ), .A(\pgld32[0] ), .B(
        \LDCHK/n3312 ), .C(\LDCHK/n3238 ), .D(\LDCHK/n3296 ) );
    snl_oai122x0 \LBUS/U594  ( .ZN(\LBUS/n_2434 ), .A(LDS), .B(\LBUS/n1448 ), 
        .C(\LBUS/ilt[0] ), .D(\LBUS/ilt[1] ), .E(\LBUS/n1449 ) );
    snl_muxi21x1 \LDIS/U164  ( .ZN(\LDIS/ldexcl[8] ), .A(\LDIS/n3135 ), .B(
        \LDIS/n3136 ), .S(\LDIS/n3134 ) );
    snl_mux21x1 \ALUSHT/U17  ( .Z(\pkdptout[4] ), .A(\ALUSHT/pkshtout[4] ), 
        .B(\ALUSHT/pkaluout[4] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U56  ( .Z(\CONS/n560 ), .A(\CONS/SACO[13] ), .B(
        \pgsdprlh[17] ) );
    snl_invx05 \SAEXE/U133  ( .ZN(\SAEXE/n426 ), .A(\SAEXE/wrd_datah ) );
    snl_invx05 \SAEXE/U97  ( .ZN(ph_tprsel_h), .A(\SAEXE/n419 ) );
    snl_ao022x1 \REGF/U497  ( .Z(\REGF/RI_PCOL[28] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[28]), .C(\stream4[28] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U520  ( .Z(\REGF/RI_PCOL[5] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[5]), .C(\stream4[5] ), .D(\REGF/n8209 ) );
    snl_ao2222x1 \REGF/U527  ( .Z(\REGF/RI_SRDA[30] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[30]), .C(\pgldi[30] ), .D(\REGF/n8210 ), .E(\stream3[30] ), .F(
        \REGF/n8211 ), .G(\pkdptout[30] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U617  ( .ZN(\REGF/RI_SPR[12] ), .A(\REGF/n8183 ), .B(
        \REGF/n8220 ), .C(\REGF/n8184 ), .D(\REGF/n8221 ), .E(\REGF/n8114 ), 
        .F(\REGF/n8218 ) );
    snl_and12x1 \REGF/U630  ( .Z(\REGF/RI_STAT[5] ), .A(\REGF/n8222 ), .B(
        PDLIN[31]) );
    snl_invx05 \MAIN/U163  ( .ZN(ph_baccwt_h), .A(\MAIN/n3615 ) );
    snl_invx05 \REGF/U787  ( .ZN(\REGF/n8134 ), .A(\pkdptout[5] ) );
    snl_invx05 \ADOSEL/U80  ( .ZN(\ADOSEL/n4088 ), .A(\pkdptout[16] ) );
    snl_xor2x0 \LDCHK/U76  ( .Z(\LDCHK/n3304 ), .A(\pgld32[17] ), .B(
        \LDCHK/pglpinff[2] ) );
    snl_nor02x1 \CONS/U38  ( .ZN(\CONS/n548 ), .A(\CONS/n549 ), .B(\CONS/n550 
        ) );
    snl_ao022x1 \MAIN/U144  ( .Z(\MAIN/ph_rrmwh ), .A(rrmw1), .B(
        \MAIN/ph_rdwr1selh ), .C(rrmw2), .D(\MAIN/ph_rdwr2selh ) );
    snl_oai112x0 \PDOSEL/U49  ( .ZN(PDLOUT[20]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n106 ), .C(\PDOSEL/n124 ), .D(\PDOSEL/n125 ) );
    snl_muxi21x1 \LDCHK/U51  ( .ZN(\LDCHK/n3246 ), .A(\LDCHK/n3271 ), .B(
        \LDCHK/n3266 ), .S(\pgld32[30] ) );
    snl_and02x1 \ALUIS/U12  ( .Z(\ALUIS/n3645 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3658 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[3]  ( .Q(\ph_segset_h[3] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[3]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_invx05 \CODEIF/U250  ( .ZN(\CODEIF/n3866 ), .A(PDLIN[0]) );
    snl_invx05 \CODEIF/U277  ( .ZN(\CODEIF/n3915 ), .A(PDLIN[16]) );
    snl_oai013x0 \LBUS/U571  ( .ZN(\LBUS/*cell*3982/U158/Z_0 ), .A(
        \LBUS/n1415 ), .B(\LBUS/n1416 ), .C(\LBUS/n1417 ), .D(\LBUS/n1418 ) );
    snl_xnor2x0 \CONS/U206  ( .ZN(\CONS/n687 ), .A(\pk_pc_h[0] ), .B(
        \pk_pcs2_h[0] ) );
    snl_and02x1 \REG_2/U157  ( .Z(\ph_cpudout[27] ), .A(\ph_segset_h[27] ), 
        .B(seg_cnfg_h) );
    snl_muxi21x1 \BLU/U411  ( .ZN(obacc), .A(\BLU/n1584 ), .B(\BLU/n1585 ), 
        .S(po_opcsel_h) );
    snl_muxi21x1 \LDIS/U181  ( .ZN(\LDIS/ldexch[29] ), .A(\LDIS/n3156 ), .B(
        \LDIS/n3155 ), .S(\LDIS/n3165 ) );
    snl_nand13x1 \LBUS/U641  ( .ZN(\LBUS/n1427 ), .A(\LBUS/temp1[2] ), .B(
        \LBUS/n1422 ), .C(\LBUS/n1603 ) );
    snl_invx05 \BLU/U390  ( .ZN(\BLU/n1470 ), .A(\pgld16[14] ) );
    snl_nand04x0 \CONS/U136  ( .ZN(\CONS/n686 ), .A(\CONS/n687 ), .B(
        \CONS/n688 ), .C(\CONS/n689 ), .D(\CONS/n690 ) );
    snl_nor02x2 \LBUS/U556  ( .ZN(up_data_lth), .A(\LBUS/n1411 ), .B(
        \LBUS/n1437 ) );
    snl_nor02x1 \LBUS/U666  ( .ZN(pgfbadrsel), .A(\LBUS/n1404 ), .B(
        \LBUS/n1452 ) );
    snl_xor2x0 \CONS/U94  ( .Z(\CONS/n612 ), .A(\pk_idcy_h[9] ), .B(
        \pk_indy_h[9] ) );
    snl_xor2x0 \CONS/U111  ( .Z(\CONS/n629 ), .A(\pk_idcw_h[6] ), .B(
        \pk_indw_h[6] ) );
    snl_xnor2x0 \CONS/U221  ( .ZN(\CONS/n705 ), .A(\pk_idcz_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_oai012x1 \BLU/U436  ( .ZN(\BLU/n1557 ), .A(\BLU/n1521 ), .B(
        \BLU/n1555 ), .C(\BLU/n1587 ) );
    snl_aoi022x1 \ALUIS/U99  ( .ZN(\ALUIS/n3694 ), .A(\stream4[2] ), .B(
        immbsel), .C(\pk_adb_h[2] ), .D(po_brsel_h) );
    snl_oai222x0 \REGF/U610  ( .ZN(\REGF/RI_SPR[19] ), .A(\REGF/n8169 ), .B(
        \REGF/n8220 ), .C(\REGF/n8170 ), .D(\REGF/n8221 ), .E(\REGF/n8093 ), 
        .F(\REGF/n8218 ) );
    snl_ffqrnx1 \CODEIF/pgfpcel_reg  ( .Q(CRCE), .D(\CODEIF/pgfpcel169 ), .RN(
        \CODEIF/n3861 ), .CP(SCLK) );
    snl_invx1 \ALUIS/U15  ( .ZN(\pgaluina[11] ), .A(\ALUIS/n3647 ) );
    snl_xor2x0 \LDCHK/U56  ( .Z(\LDCHK/n3256 ), .A(\LDCHK/n3278 ), .B(
        \LDCHK/n3279 ) );
    snl_oai022x1 \REGF/U637  ( .ZN(\REGF/RI_TBAI[21] ), .A(\REGF/n8225 ), .B(
        \REGF/n8155 ), .C(\REGF/n8226 ), .D(\REGF/n8156 ) );
    snl_invx05 \REGF/U780  ( .ZN(\REGF/n8207 ), .A(\pgregadrh[0] ) );
    snl_nand02x1 \ADOSEL/U87  ( .ZN(\ADOSEL/n4100 ), .A(\pgbluext[3] ), .B(
        \ADOSEL/n4156 ) );
    snl_ao012x1 \MAIN/U143  ( .Z(ph_aluovf_h), .A(wacc), .B(pkaluovf), .C(
        \MAIN/accovf ) );
    snl_and02x1 \MAIN/U164  ( .Z(\MAIN/excep_valid ), .A(pk_excp_h), .B(
        \MAIN/excep_enable ) );
    snl_xor2x0 \LDCHK/U71  ( .Z(\LDCHK/n3300 ), .A(\pgld32[14] ), .B(
        \pgld32[15] ) );
    snl_oai112x0 \PDOSEL/U69  ( .ZN(PDLOUT[18]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n104 ), .C(\PDOSEL/n160 ), .D(\PDOSEL/n161 ) );
    snl_ao022x1 \REGF/U507  ( .Z(\REGF/RI_PCOL[18] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[18]), .C(\stream4[18] ), .D(\REGF/n8209 ) );
    snl_invx05 \REGF/U742  ( .ZN(\REGF/n8091 ), .A(\pgldi[19] ) );
    snl_invx05 \ADOSEL/U45  ( .ZN(\ADOSEL/n4116 ), .A(\pkdptout[25] ) );
    snl_invx05 \CODEIF/U257  ( .ZN(\CODEIF/n3891 ), .A(PDLIN[8]) );
    snl_nand02x1 \ALUIS/U32  ( .ZN(\pgaluina[16] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3674 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[1]  ( .Q(\ph_segset_h[1] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[1]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_xnor2x0 \CONS/U226  ( .ZN(\CONS/n709 ), .A(\pk_idcz_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \BLU/U431  ( .ZN(oltff), .A(\BLU/n1518 ) );
    snl_invx05 \CODEIF/U270  ( .ZN(\CODEIF/n3869 ), .A(\CODEIF/pfctr[1] ) );
    snl_muxi21x1 \LDIS/U186  ( .ZN(\LDIS/ldexch[24] ), .A(\LDIS/n3136 ), .B(
        \LDIS/n3135 ), .S(\LDIS/n3165 ) );
    snl_invx05 \LBUS/U661  ( .ZN(\LBUS/*cell*3982/U71/CONTROL1 ), .A(
        \LBUS/n1401 ) );
    snl_xor2x0 \CONS/U116  ( .Z(\CONS/n634 ), .A(\pk_idcw_h[18] ), .B(
        \pk_indw_h[18] ) );
    snl_xor2x0 \CONS/U93  ( .Z(\CONS/n611 ), .A(\pk_idcy_h[4] ), .B(
        \pk_indy_h[4] ) );
    snl_aoi122x0 \LBUS/U646  ( .ZN(\LBUS/n1400 ), .A(\LBUS/n1435 ), .B(
        \LBUS/n1436 ), .C(\LBUS/n1590 ), .D(word32odtrh), .E(ph_lberr) );
    snl_nand03x0 \CONS/U131  ( .ZN(\CONS/n563 ), .A(\CONS/n671 ), .B(
        \CONS/n672 ), .C(\CONS/n673 ) );
    snl_xnor2x0 \CONS/U201  ( .ZN(\CONS/n683 ), .A(\pk_pc_h[11] ), .B(
        \pk_pcs2_h[11] ) );
    snl_and02x1 \REG_2/U150  ( .Z(\ph_cpudout[20] ), .A(\ph_segset_h[20] ), 
        .B(seg_cnfg_h) );
    snl_nand02x1 \BLU/U397  ( .ZN(\BLU/n1477 ), .A(\BLU/n1565 ), .B(
        \BLU/n1562 ) );
    snl_oa2222x1 \BLU/U416  ( .Z(\BLU/n1513 ), .A(\BLU/n1474 ), .B(\BLU/n1476 
        ), .C(\BLU/n1471 ), .D(\BLU/n1473 ), .E(\BLU/n1468 ), .F(\BLU/n1470 ), 
        .G(\BLU/n1465 ), .H(\BLU/n1467 ) );
    snl_nand02x2 \ALUIS/U7  ( .ZN(\pgaluina[12] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3670 ) );
    snl_or03x1 \LBUS/U576  ( .Z(\LBUS/nlt[5] ), .A(ph_d53lth), .B(ph_d20lth), 
        .C(\LBUS/n1434 ) );
    snl_nand12x1 \LBUS/U628  ( .ZN(\LBUS/n1445 ), .A(\LBUS/n1597 ), .B(
        \LBUS/n1596 ) );
    snl_nand02x1 \PDOSEL/U153  ( .ZN(\PDOSEL/n130 ), .A(CDIN[19]), .B(
        \PDOSEL/n119 ) );
    snl_oai012x1 \LDCHK/U94  ( .ZN(\LDCHK/n3237 ), .A(\LDCHK/n3247 ), .B(
        \LDCHK/n3250 ), .C(ph_pdlen_h) );
    snl_invx05 \REGF/U800  ( .ZN(\REGF/n8083 ), .A(\pkdptout[22] ) );
    snl_oai122x0 \CODEIF/U239  ( .ZN(\CODEIF/pfctr415[18] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3920 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3921 ), .E(
        \CODEIF/n3922 ) );
    snl_xnor2x0 \CONS/U248  ( .ZN(\CONS/n732 ), .A(\pk_idcx_h[20] ), .B(
        \pk_indx_h[20] ) );
    snl_mux21x1 \SHTCD/U14  ( .Z(\phshtd[2] ), .A(\pgld16[2] ), .B(
        \stream4[2] ), .S(immbsel) );
    snl_or04x1 \REGF/U659  ( .Z(\REGF/RO_PSTA[17] ), .A(\REGF/RO_EST2[2] ), 
        .B(\REGF/RO_EST2[1] ), .C(\REGF/RO_EST2[15] ), .D(\REGF/RO_EST2[0] )
         );
    snl_invx05 \REGF/U765  ( .ZN(\REGF/n8166 ), .A(\pgsdprlh[21] ) );
    snl_invx05 \REGF/U827  ( .ZN(\REGF/n8224 ), .A(\REGF/n8232 ) );
    snl_invx05 \ADOSEL/U62  ( .ZN(\ADOSEL/n4135 ), .A(\pkdptout[15] ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[0]  ( .Q(CA[0]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3765 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_xnor2x0 \CONS/U178  ( .ZN(\CONS/n663 ), .A(\pgsdprlh[19] ), .B(
        \pk_saco_lh[19] ) );
    snl_muxi21x1 \LDIS/U163  ( .ZN(\LDIS/ldexcl[9] ), .A(\LDIS/n3132 ), .B(
        \LDIS/n3133 ), .S(\LDIS/n3134 ) );
    snl_nor03x4 \ALUSHT/U10  ( .ZN(\ALUSHT/n3112 ), .A(\poshtfnc[2] ), .B(
        \poshtfnc[1] ), .C(\poshtfnc[0] ) );
    snl_xor2x0 \CONS/U51  ( .Z(\CONS/n573 ), .A(\pk_saco_lh[15] ), .B(
        \pgsdprlh[15] ) );
    snl_and02x1 \SAEXE/U134  ( .Z(\SAEXE/sequen ), .A(\pk_psae_h[6] ), .B(
        \SAEXE/n429 ) );
    snl_aoi012x1 \LBUS/U593  ( .ZN(\LBUS/ldoe966 ), .A(ph_lbwrh), .B(
        \LBUS/nlt[3] ), .C(\LBUS/n1399 ) );
    snl_oai2222x0 \REGF/U363  ( .ZN(\REGF/RI_SRA12M[8] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8126 ), .C(\REGF/n8124 ), .D(\REGF/n8051 ), .E(\REGF/n8191 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8192 ) );
    snl_invx2 \REGF/U378  ( .ZN(\REGF/n8059 ), .A(\ph_pdis_h[1] ) );
    snl_and02x1 \REGF/U569  ( .Z(\REGF/RO_LPSAS2156[11] ), .A(
        \REGF/RO_PSASH[15] ), .B(ph_sastlth) );
    snl_xnor2x0 \LDCHK/U110  ( .ZN(\LDCHK/n3287 ), .A(\pgmuxout[12] ), .B(
        \pgmuxout[10] ) );
    snl_ao2222x1 \REGF/U555  ( .Z(\REGF/RI_SRDA[2] ), .A(PDLIN[2]), .B(
        \ph_pdis_h[9] ), .C(\pgldi[2] ), .D(\REGF/n8210 ), .E(\stream3[2] ), 
        .F(\REGF/n8211 ), .G(\pkdptout[2] ), .H(\REGF/n8212 ) );
    snl_invx05 \REGF/U665  ( .ZN(\REGF/n8117 ), .A(PDLIN[11]) );
    snl_ao222x1 \CODEIF/U199  ( .Z(\CODEIF/n3846 ), .A(PA[8]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[5] ), .E(cif_byte), .F(PDLIN[5])
         );
    snl_xor2x0 \CODEIF/U295  ( .Z(\CODEIF/n3957 ), .A(\CODEIF/n3958 ), .B(CDIN
        [0]) );
    snl_xor2x0 \CODEIF/U305  ( .Z(\CODEIF/n3950 ), .A(\CODEIF/n3972 ), .B(
        \CODEIF/n3973 ) );
    snl_aoi022x1 \ALUIS/U135  ( .ZN(\ALUIS/n3716 ), .A(\stream4[13] ), .B(
        immbsel), .C(\pk_adb_h[13] ), .D(po_brsel_h) );
    snl_invx05 \BLU/U372  ( .ZN(\BLU/n1494 ), .A(\pgld16[6] ) );
    snl_xor2x0 \CODEIF/U322  ( .Z(\CODEIF/n3999 ), .A(CDOUT[51]), .B(CDOUT[47]
        ) );
    snl_aoi012x1 \ALUIS/U112  ( .ZN(\ALUIS/n3737 ), .A(\pgldi[23] ), .B(
        srcbsel), .C(allfbsel) );
    snl_nor02x1 \BLU/U355  ( .ZN(\BLU/n1570 ), .A(\BLU/n1564 ), .B(
        \pgbitnoh[1] ) );
    snl_xor2x0 \LDCHK/U38  ( .Z(\LDCHK/n3247 ), .A(\LDCHK/n3248 ), .B(
        \LDCHK/n3249 ) );
    snl_oai012x1 \LDIS/U144  ( .ZN(\pgldi[30] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3130 ), .C(\LDIS/n3115 ) );
    snl_mux21x1 \ALUSHT/U37  ( .Z(\pkdptout[15] ), .A(\ALUSHT/pkshtout[15] ), 
        .B(\ALUSHT/pkaluout[15] ), .S(\ALUSHT/n3112 ) );
    snl_nand02x1 \LBUS/U684  ( .ZN(\LBUS/n1440 ), .A(\LBUS/n1460 ), .B(
        \LBUS/ilt[1] ) );
    snl_oai013x0 \SAEXE/U113  ( .ZN(phadrinch), .A(\SAEXE/n424 ), .B(
        \pk_psae_h[3] ), .C(\SAEXE/n413 ), .D(\SAEXE/n415 ) );
    snl_xor2x0 \CONS/U76  ( .Z(\CONS/n594 ), .A(\pk_pcs1_h[10] ), .B(
        \pk_pc_h[10] ) );
    snl_oai012x1 \PDOSEL/U20  ( .ZN(PDH[36]), .A(\PDOSEL/n80 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nor03x0 \MAIN/U136  ( .ZN(\MAIN/single_write ), .A(\MAIN/n3630 ), .B(
        pkaccovf), .C(pgadrovfh) );
    snl_nand02x1 \ADOSEL/U106  ( .ZN(\ADOSEL/n4136 ), .A(\pgbluext[31] ), .B(
        \ADOSEL/n4156 ) );
    snl_and03x1 \SAEXE/U108  ( .Z(phbnolth), .A(\SAEXE/bnolth ), .B(ph_bitsrch
        ), .C(\SAEXE/stage_1st ) );
    snl_nand02x1 \CODEIF/U339  ( .ZN(\CODEIF/n3895 ), .A(\CODEIF/n3945 ), .B(
        \CODEIF/pgctrinc[9] ) );
    snl_nand02x1 \ALUIS/U60  ( .ZN(\pgaluinb[12] ), .A(\ALUIS/n3714 ), .B(
        \ALUIS/n3715 ) );
    snl_aoi022x1 \ALUIS/U109  ( .ZN(\ALUIS/n3740 ), .A(\stream4[25] ), .B(
        immbsel), .C(\pk_adb_h[25] ), .D(po_brsel_h) );
    snl_oai222x0 \REGF/U572  ( .ZN(\REGF/RI_ACC[29] ), .A(\REGF/n8063 ), .B(
        \REGF/n8215 ), .C(\REGF/n8064 ), .D(\REGF/n8216 ), .E(\REGF/n8155 ), 
        .F(\REGF/n8217 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[9]  ( .Q(CA[9]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3861 ), .SD(\CODEIF/n3850 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_nand02x1 \ALUIS/U47  ( .ZN(\pgaluina[31] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3689 ) );
    snl_and02x1 \UPIF/U15  ( .Z(\ph_pdis_h[2] ), .A(\pk_rread_h[61] ), .B(
        \UPIF/n1046 ) );
    snl_invx05 \BLU/U369  ( .ZN(\BLU/n1491 ), .A(\pgld16[7] ) );
    snl_oai012x2 \REGF/U386  ( .ZN(\REGF/n8229 ), .A(ph_srcadr2_h), .B(
        ph_srcadr1_h), .C(\REGF/n8228 ) );
    snl_oai022x1 \REGF/U469  ( .ZN(\REGF/RI_DPR[24] ), .A(\REGF/n8157 ), .B(
        \REGF/n8151 ), .C(\REGF/n8152 ), .D(\REGF/n8158 ) );
    snl_oai022x1 \REGF/U642  ( .ZN(\REGF/RI_TBAI[15] ), .A(\REGF/n8225 ), .B(
        \REGF/n8093 ), .C(\REGF/n8226 ), .D(\REGF/n8169 ) );
    snl_muxi21x1 \LDIS/U178  ( .ZN(\LDIS/ldexcl[0] ), .A(\LDIS/n3163 ), .B(
        \LDIS/n3164 ), .S(\LDIS/n3134 ) );
    snl_invx05 \LBUS/U588  ( .ZN(LDS), .A(\LBUS/temp[3] ) );
    snl_invx05 \ADOSEL/U79  ( .ZN(\ADOSEL/n4090 ), .A(\pkdptout[0] ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[6]  ( .Q(\CODEIF/pfctr[6] ), .D(
        \CODEIF/pfctr415[6] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nor03x0 \LBUS/U614  ( .ZN(\LBUS/n1590 ), .A(\LBUS/n1452 ), .B(
        \LBUS/ilt[5] ), .C(\LBUS/n1463 ) );
    snl_oai122x0 \CODEIF/U222  ( .ZN(\CODEIF/pfctr415[1] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3869 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3870 ), .E(
        \CODEIF/n3871 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[15]  ( .Q(\CODEIF/pfctr[15] ), .D(
        \CODEIF/pfctr415[15] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_invx05 \CONS/U163  ( .ZN(\CONS/n650 ), .A(\CONS/n552 ) );
    snl_xnor2x0 \CONS/U253  ( .ZN(\CONS/n735 ), .A(\pk_idcx_h[14] ), .B(
        \pk_indx_h[14] ) );
    snl_muxi21x1 \BLU/U444  ( .ZN(\BLU/n1584 ), .A(\BLU/n1583 ), .B(
        \BLU/n1582 ), .S(po_cmfsel_h) );
    snl_invx05 \REGF/U759  ( .ZN(\REGF/n8202 ), .A(\pgsdprlh[3] ) );
    snl_ao222x1 \CODEIF/U205  ( .Z(\CODEIF/n3852 ), .A(PA[14]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[11] ), .E(cif_byte), .F(PDLIN[11]
        ) );
    snl_xnor2x0 \CODEIF/U395  ( .ZN(\CODEIF/n3990 ), .A(CDIN[7]), .B(CDIN[8])
         );
    snl_xnor2x0 \CODEIF/U414  ( .ZN(\CODEIF/n4010 ), .A(CDOUT[29]), .B(CDOUT
        [25]) );
    snl_sffqenrnx1 \CODEIF/fm_config_reg[1]  ( .Q(\CODEIF/fm_config[1] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEIF/n3862 ), .SD(PDLIN[1]), .SE(cnfg_write_h
        ), .CP(SCLK) );
    snl_xnor2x0 \CONS/U274  ( .ZN(\CONS/n338 ), .A(\pk_idcw_h[10] ), .B(
        \pk_indw_h[10] ) );
    snl_invx05 \LBUS/U633  ( .ZN(\LBUS/n1459 ), .A(\LBUS/ph_lbusylth ) );
    snl_nor03x0 \CONS/U144  ( .ZN(\CONS/n531 ), .A(\CONS/n606 ), .B(
        \CONS/n604 ), .C(\CONS/n605 ) );
    snl_nand02x1 \PDOSEL/U148  ( .ZN(\PDOSEL/n154 ), .A(CDIN[22]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \PDOSEL/U97  ( .ZN(\PDOSEL/n103 ), .A(CDIN[49]) );
    snl_ao022x1 \REGF/U407  ( .Z(\REGF/RI_PCOH[26] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[26]), .C(\stream4[58] ), .D(\REGF/n8053 ) );
    snl_ao022x1 \REGF/U420  ( .Z(\REGF/RI_PCOH[13] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[13]), .C(\stream4[45] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U597  ( .ZN(\REGF/RI_ACC[4] ), .A(\REGF/n8136 ), .B(
        \REGF/n8215 ), .C(\REGF/n8137 ), .D(\REGF/n8216 ), .E(\REGF/n8138 ), 
        .F(\REGF/n8217 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[8]  ( .Q(\ph_segset_h[8] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[8]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_invx05 \REGF/U680  ( .ZN(\REGF/n8156 ), .A(\pgsdprhh[29] ) );
    snl_invx05 \REGF/U737  ( .ZN(\REGF/n8079 ), .A(\pgldi[23] ) );
    snl_oai122x0 \ADOSEL/U30  ( .ZN(\pgmuxout[19] ), .A(\ADOSEL/n4099 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4098 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4142 ) );
    snl_nor02x1 \PDOSEL/U126  ( .ZN(\PDOSEL/n153 ), .A(\pk_pdo_h[17] ), .B(
        \ph_cpudout[17] ) );
    snl_xor2x0 \CONS/U88  ( .Z(\CONS/n606 ), .A(\pk_idcz_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_invx05 \REGF/U710  ( .ZN(\REGF/n8147 ), .A(PDLIN[1]) );
    snl_oai122x0 \ADOSEL/U17  ( .ZN(\pgmuxout[6] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4107 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4108 ), .E(
        \ADOSEL/n4109 ) );
    snl_invx05 \PDOSEL/U101  ( .ZN(\PDOSEL/n99 ), .A(CDIN[45]) );
    snl_oai222x0 \REGF/U619  ( .ZN(\REGF/RI_SPR[10] ), .A(\REGF/n8187 ), .B(
        \REGF/n8220 ), .C(\REGF/n8188 ), .D(\REGF/n8221 ), .E(\REGF/n8120 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U789  ( .ZN(\REGF/n8140 ), .A(\pkdptout[3] ) );
    snl_nand02x1 \CODEIF/U357  ( .ZN(\CODEIF/n3868 ), .A(\CODEIF/pgctrinc[0] ), 
        .B(\CODEIF/n3945 ) );
    snl_nand02x1 \CODEIF/U370  ( .ZN(\CODEIF/n3962 ), .A(write_pr_h), .B(
        \CODEIF/write_prtect ) );
    snl_nand02x2 \ALUIS/U29  ( .ZN(\pgaluina[15] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3673 ) );
    snl_aoi022x1 \ALUIS/U85  ( .ZN(\ALUIS/n3704 ), .A(\stream4[7] ), .B(
        immbsel), .C(\pk_adb_h[7] ), .D(po_brsel_h) );
    snl_aoi012x1 \ALUIS/U140  ( .ZN(\ALUIS/n3711 ), .A(\pgldi[10] ), .B(
        srcbsel), .C(allfbsel) );
    snl_oai022x1 \BLU/U307  ( .ZN(\pkbludgh[9] ), .A(\BLU/n1464 ), .B(
        \BLU/n1483 ), .C(\BLU/n1484 ), .D(\BLU/n1485 ) );
    snl_nand02x1 \ALUIS/U167  ( .ZN(\ALUIS/n3675 ), .A(\pk_ada_h[17] ), .B(
        po_arsel_h) );
    snl_ao022x1 \BLUOS/U17  ( .Z(\pgbluext[29] ), .A(\pkbludgh[13] ), .B(
        ph_bit_h), .C(\pkdptout[13] ), .D(ph_word16_h) );
    snl_invx05 \MAIN/U158  ( .ZN(\MAIN/*cell*4603/U7/CONTROL1 ), .A(
        \MAIN/n3617 ) );
    snl_ao022x1 \LDIS/U116  ( .Z(\pgldi[9] ), .A(\pgld32[9] ), .B(ph_word32_h), 
        .C(\pgld16[9] ), .D(ph_word16_h) );
    snl_invx05 \LDIS/U226  ( .ZN(\LDIS/n3152 ), .A(LIN[31]) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[0]  ( .Q(\REG_2/RETCNT[0] ), .D(
        \REG_2/ph_retcnt_h[0] ), .EN(\REG_2/n517 ), .RN(\REG_2/n436 ), .SD(
        \REG_2/ncnt1[0] ), .SE(ph_d20lth), .CP(SCLK) );
    snl_oai012x1 \LDIS/U131  ( .ZN(\pgldi[17] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3117 ), .C(\LDIS/n3115 ) );
    snl_ao022x1 \CMPX/U20  ( .Z(ph_wrdsrc_h), .A(ph_wrdsrch), .B(ph_saexe_sth), 
        .C(po_wrdsrc_h), .D(\CMPX/n1047 ) );
    snl_oai112x0 \PDOSEL/U72  ( .ZN(PDLOUT[23]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n109 ), .C(\PDOSEL/n164 ), .D(\PDOSEL/n177 ) );
    snl_nand02x1 \SAEXE/U141  ( .ZN(\SAEXE/n420 ), .A(\SAEXE/srcwrit ), .B(
        ph_saexe_sth) );
    snl_mux21x1 \ALUSHT/U42  ( .Z(\pkdptout[10] ), .A(\ALUSHT/pkshtout[10] ), 
        .B(\ALUSHT/pkaluout[10] ), .S(\ALUSHT/n3112 ) );
    snl_xnor2x0 \CONS/U186  ( .ZN(\CONS/n666 ), .A(\pk_saco_lh[2] ), .B(
        \pgsdprlh[2] ) );
    snl_oai112x0 \PDOSEL/U55  ( .ZN(PDLOUT[27]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n113 ), .C(\PDOSEL/n134 ), .D(\PDOSEL/n135 ) );
    snl_xor2x0 \CODEIF/U362  ( .Z(\CODEIF/n3937 ), .A(CDOUT[45]), .B(
        \CODEIF/n4022 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[15]  ( .Q(CA[15]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3856 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_aoi022x1 \BLU/U320  ( .ZN(\BLU/n1521 ), .A(\BLU/n1522 ), .B(
        \BLU/n1523 ), .C(\BLU/n1524 ), .D(\BLU/n1525 ) );
    snl_nand02x1 \ALUIS/U152  ( .ZN(\ALUIS/n3688 ), .A(\pk_ada_h[30] ), .B(
        po_arsel_h) );
    snl_ffqx1 \MAIN/LBAOVFH_reg  ( .Q(\MAIN/LBAOVFH ), .D(ph_lbaovf), .CP(SCLK
        ) );
    snl_invx05 \LDIS/U201  ( .ZN(\LDIS/n3145 ), .A(LIN[3]) );
    snl_invx2 \SAEXE/U99  ( .ZN(ph_dregsl_h), .A(\SAEXE/n420 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[18]  ( .Q(\CODEIF/pfctr[18] ), .D(
        \CODEIF/pfctr415[18] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nor02x1 \CMPX/U15  ( .ZN(\CMPX/n1049 ), .A(phadrinch), .B(\CMPX/n1047 
        ) );
    snl_oai112x0 \PDOSEL/U60  ( .ZN(PDLOUT[2]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n78 ), .C(\PDOSEL/n144 ), .D(\PDOSEL/n145 ) );
    snl_oai022x1 \BLU/U315  ( .ZN(\pkbludgh[1] ), .A(\BLU/n1464 ), .B(
        \BLU/n1507 ), .C(\BLU/n1508 ), .D(\BLU/n1509 ) );
    snl_ao022x1 \BLUOS/U22  ( .Z(\pgbluext[3] ), .A(\pkbludgh[3] ), .B(
        ph_bit_h), .C(\pkdptout[3] ), .D(ph_word16_h) );
    snl_ao022x1 \LDIS/U104  ( .Z(\pgldi[3] ), .A(ph_word32_h), .B(\pgld32[3] ), 
        .C(\pgld16[3] ), .D(ph_word16_h) );
    snl_nor02x1 \CONS/U36  ( .ZN(\CONS/n545 ), .A(\CONS/n543 ), .B(\CONS/n546 
        ) );
    snl_xor2x0 \LDCHK/U78  ( .Z(\LDCHK/n3305 ), .A(\LDCHK/pglpinff[3] ), .B(
        \pgld32[28] ) );
    snl_ao022x1 \LDIS/U123  ( .Z(\pgld16[12] ), .A(ph_selldl), .B(\pgld32[12] 
        ), .C(ph_selldh), .D(\pgld32[28] ) );
    snl_xnor2x0 \CONS/U194  ( .ZN(\CONS/n680 ), .A(\pk_pc_h[17] ), .B(
        \pk_pcs2_h[17] ) );
    snl_oai112x0 \PDOSEL/U47  ( .ZN(PDLOUT[1]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n77 ), .C(\PDOSEL/n120 ), .D(\PDOSEL/n121 ) );
    snl_nand02x3 \REGF/U394  ( .ZN(\REGF/n8056 ), .A(ph_rgfile_h), .B(
        \REGF/n8059 ) );
    snl_ao2222x1 \REGF/U529  ( .Z(\REGF/RI_SRDA[28] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[28]), .C(\pgldi[28] ), .D(\REGF/n8210 ), .E(\stream3[28] ), .F(
        \REGF/n8211 ), .G(\pkdptout[28] ), .H(\REGF/n8212 ) );
    snl_nand02x1 \CODEIF/U345  ( .ZN(\CODEIF/n3877 ), .A(\CODEIF/pgctrinc[3] ), 
        .B(\CODEIF/n3945 ) );
    snl_nand02x1 \ALUIS/U175  ( .ZN(\ALUIS/n3658 ), .A(\pk_ada_h[0] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U213  ( .ZN(\LDIS/n3132 ), .A(LIN[9]) );
    snl_nor02x1 \BLU/U332  ( .ZN(\BLU/n1469 ), .A(\BLU/n1546 ), .B(\BLU/n1547 
        ) );
    snl_oai222x0 \REGF/U585  ( .ZN(\REGF/RI_ACC[16] ), .A(\REGF/n8100 ), .B(
        \REGF/n8215 ), .C(\REGF/n8101 ), .D(\REGF/n8216 ), .E(\REGF/n8102 ), 
        .F(\REGF/n8217 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[4]  ( .Q(CA[4]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3845 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_ffqrnx1 \MAIN/cstregw_tap1_reg  ( .Q(\MAIN/cstregw_tap1 ), .D(
        \MAIN/*cell*4603/U10/CONTROL1 ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_ao022x1 \REGF/U415  ( .Z(\REGF/RI_PCOH[18] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[18]), .C(\stream4[50] ), .D(\REGF/n8053 ) );
    snl_ao022x1 \REGF/U432  ( .Z(\REGF/RI_PCOH[1] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[1]), .C(\stream4[33] ), .D(\REGF/n8053 ) );
    snl_invx05 \REGF/U692  ( .ZN(\REGF/n8167 ), .A(\pgregadrh[20] ) );
    snl_invx05 \REGF/U702  ( .ZN(\REGF/n8177 ), .A(\pgregadrh[15] ) );
    snl_invx05 \REGF/U725  ( .ZN(\REGF/n8142 ), .A(\pgldi[2] ) );
    snl_invx05 \CODEIF/U279  ( .ZN(\CODEIF/n3912 ), .A(PDLIN[15]) );
    snl_xnor2x0 \CONS/U208  ( .ZN(\CONS/n697 ), .A(\pk_pc_h[4] ), .B(
        \pk_pcs1_h[4] ) );
    snl_and02x1 \REG_2/U159  ( .Z(\ph_cpudout[29] ), .A(\ph_segset_h[29] ), 
        .B(seg_cnfg_h) );
    snl_oai122x0 \ADOSEL/U22  ( .ZN(\pgmuxout[11] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4122 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4123 ), .E(
        \ADOSEL/n4124 ) );
    snl_nor03x0 \CONS/U138  ( .ZN(\CONS/n691 ), .A(\CONS/n593 ), .B(
        \CONS/n591 ), .C(\CONS/n592 ) );
    snl_aoi112x0 \PDOSEL/U134  ( .ZN(\PDOSEL/n179 ), .A(\pgfdout[0] ), .B(
        \PDOSEL/n226 ), .C(\pk_pdo_h[0] ), .D(\ph_cpudout[0] ) );
    snl_ffqsnx1 \LBUS/ldoe_reg  ( .Q(LCNT), .D(\LBUS/ldoe966 ), .SN(n10734), 
        .CP(SCLK) );
    snl_invx05 \LBUS/U668  ( .ZN(\LBUS/n1437 ), .A(ph_lpdilth) );
    snl_nor02x1 \PDOSEL/U113  ( .ZN(\PDOSEL/n129 ), .A(\ph_cpudout[3] ), .B(
        \pk_pdo_h[3] ) );
    snl_nand02x1 \LBUS/U558  ( .ZN(phrstith), .A(ph_lbwrh), .B(\LBUS/temp1[2] 
        ) );
    snl_invx05 \REGF/U809  ( .ZN(\REGF/n8107 ), .A(\pkdptout[14] ) );
    snl_oai122x0 \CODEIF/U230  ( .ZN(\CODEIF/pfctr415[9] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3893 ), .C(\CODEIF/n3894 ), .D(\CODEIF/n3867 ), .E(
        \CODEIF/n3895 ) );
    snl_xnor2x0 \CODEIF/U421  ( .ZN(\CODEIF/n4043 ), .A(CDOUT[12]), .B(CDOUT
        [7]) );
    snl_aoi022x1 \ALUIS/U97  ( .ZN(\ALUIS/n3750 ), .A(\stream4[30] ), .B(
        immbsel), .C(\pk_adb_h[30] ), .D(po_brsel_h) );
    snl_mux21x1 \BLU/U438  ( .Z(\BLU/n1554 ), .A(\BLU/n1574 ), .B(
        \pk_stat_h[1] ), .S(eaccbsel) );
    snl_sffqenrnx1 \LDCHK/pglpinff_reg[2]  ( .Q(\LDCHK/pglpinff[2] ), .D(1'b0), 
        .EN(1'b1), .RN(n10733), .SD(\LDCHK/lpex[2] ), .SE(ph_lpdilth), .CP(
        SCLK) );
    snl_nand03x0 \LBUS/U606  ( .ZN(\LBUS/n1416 ), .A(\LBUS/n1458 ), .B(
        \LBUS/n1425 ), .C(\LBUS/n1459 ) );
    snl_xnor2x0 \CONS/U171  ( .ZN(\CONS/n553 ), .A(\pk_saco_hh[28] ), .B(
        \pgsdprhh[28] ) );
    snl_xnor2x0 \CONS/U241  ( .ZN(\CONS/n721 ), .A(\pk_idcy_h[13] ), .B(
        \pk_indy_h[13] ) );
    snl_nor02x2 \CODEIF/U217  ( .ZN(\CODEIF/n3945 ), .A(\CODEIF/n3944 ), .B(
        cnt_write_h) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[18]  ( .Q(CA[18]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3859 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_sffqrnx1 \MAIN/POL_STH_reg  ( .Q(\MAIN/POL_STH ), .D(pol_status), .RN(
        \MAIN/n3611 ), .SD(1'b0), .SE(\MAIN/sw_end ), .CP(SCLK) );
    snl_xnor2x0 \CONS/U266  ( .ZN(\CONS/n741 ), .A(\pk_idcw_h[1] ), .B(
        \pk_indw_h[1] ) );
    snl_ao022x1 \REG_2/U137  ( .Z(\ph_cpudout[7] ), .A(\ph_segset_h[7] ), .B(
        seg_cnfg_h), .C(ret_cont_h), .D(\REG_2/ph_retcnt_h[7] ) );
    snl_xnor2x0 \CODEIF/U387  ( .ZN(\CODEIF/n3983 ), .A(CDIN[20]), .B(CPIN[1])
         );
    snl_xor2x0 \CODEIF/U406  ( .Z(\CODEIF/n3936 ), .A(\CODEIF/n4000 ), .B(
        \CODEIF/n4038 ) );
    snl_invx05 \LBUS/U621  ( .ZN(\LBUS/n1439 ), .A(stage_b) );
    snl_invx2 U9 ( .ZN(n10736), .A(n10737) );
    snl_oai2222x0 \REGF/U356  ( .ZN(\REGF/RI_SRA12M[19] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8093 ), .C(\REGF/n8091 ), .D(\REGF/n8051 ), .E(\REGF/n8169 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8170 ) );
    snl_ao2222x1 \REGF/U547  ( .Z(\REGF/RI_SRDA[10] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[10]), .C(\pgldi[10] ), .D(\REGF/n8210 ), .E(\stream3[10] ), .F(
        \REGF/n8211 ), .G(\pkdptout[10] ), .H(\REGF/n8212 ) );
    snl_invx05 \REGF/U677  ( .ZN(\REGF/n8058 ), .A(PDLIN[31]) );
    snl_nand12x1 \MAIN/U124  ( .ZN(\MAIN/*cell*4603/U15/CONTROL1 ), .A(
        \MAIN/*cell*4603/U1/CONTROL1 ), .B(\MAIN/n3616 ) );
    snl_nand03x0 \CONS/U156  ( .ZN(\CONS/n734 ), .A(\CONS/n735 ), .B(
        \CONS/n736 ), .C(\CONS/n737 ) );
    snl_invx05 \PDOSEL/U85  ( .ZN(\PDOSEL/n78 ), .A(CDIN[34]) );
    snl_nor02x1 \LDCHK/U31  ( .ZN(LPOUT[0]), .A(\LDCHK/n3231 ), .B(
        \LDCHK/n3232 ) );
    snl_oai012x1 \PDOSEL/U29  ( .ZN(PDH[45]), .A(\PDOSEL/n99 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nand02x1 \ALUIS/U72  ( .ZN(\pgaluinb[24] ), .A(\ALUIS/n3738 ), .B(
        \ALUIS/n3739 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[5]  ( .Q(\ph_segset_h[5] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[5]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_oai022x1 \REGF/U371  ( .ZN(\REGF/RI_TBAI[19] ), .A(\REGF/n8225 ), .B(
        \REGF/n8081 ), .C(\REGF/n8226 ), .D(\REGF/n8159 ) );
    snl_nand02x1 \ALUIS/U55  ( .ZN(\pgaluinb[7] ), .A(\ALUIS/n3704 ), .B(
        \ALUIS/n3705 ) );
    snl_xnor2x0 \LDCHK/U119  ( .ZN(\LDCHK/n3313 ), .A(\pgld32[8] ), .B(
        \pgld32[11] ) );
    snl_oai2222x1 \REGF/U387  ( .ZN(\REGF/RI_SRA12M[23] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8081 ), .C(\REGF/n8079 ), .D(\REGF/n8051 ), .E(\REGF/n8159 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8161 ) );
    snl_ao022x1 \REGF/U406  ( .Z(\REGF/RI_PCOH[27] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[27]), .C(\stream4[59] ), .D(\REGF/n8053 ) );
    snl_ao022x1 \REGF/U429  ( .Z(\REGF/RI_PCOH[4] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[4]), .C(\stream4[36] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U447  ( .ZN(\REGF/RI_EACC[18] ), .A(\REGF/n8094 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8095 ), .E(\REGF/n8096 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U460  ( .ZN(\REGF/RI_EACC[5] ), .A(\REGF/n8133 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8134 ), .E(\REGF/n8135 ), 
        .F(\REGF/n8059 ) );
    snl_and02x1 \REGF/U560  ( .Z(\REGF/RO_LPSAS2156[2] ), .A(ph_sastlth), .B(
        \REGF/RO_EST1[4] ) );
    snl_oai022x1 \REGF/U650  ( .ZN(\REGF/RI_TBAI[4] ), .A(\REGF/n8225 ), .B(
        \REGF/n8126 ), .C(\REGF/n8226 ), .D(\REGF/n8191 ) );
    snl_invx05 \REGF/U750  ( .ZN(\REGF/n8115 ), .A(\pgldi[11] ) );
    snl_sffqenrnx1 \REGF/IRO_STAT1_reg  ( .Q(\REGF/RO_DDCS[25] ), .D(
        \pk_stat_h[1] ), .EN(\REGF/n8269 ), .RN(\REGF/n8052 ), .SD(1'b0), .SE(
        \pk_rwrit_h[44] ), .CP(SCLK) );
    snl_mux21x1 \ALUSHT/U19  ( .Z(\pkdptout[31] ), .A(\ALUSHT/pkshtout[31] ), 
        .B(\ALUSHT/pkaluout[31] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U58  ( .Z(\CONS/n562 ), .A(\CONS/SACO[7] ), .B(
        \pgsdprlh[11] ) );
    snl_invx05 \CONS/U43  ( .ZN(\CONS/n540 ), .A(ph_lwdsrc_h) );
    snl_invx05 \SAEXE/U126  ( .ZN(\SAEXE/n428 ), .A(\SAEXE/stage_1st ) );
    snl_invx05 \ADOSEL/U57  ( .ZN(\ADOSEL/n4102 ), .A(\pkdptout[4] ) );
    snl_invx05 \CODEIF/U287  ( .ZN(\CODEIF/n3900 ), .A(PDLIN[11]) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[11]  ( .Q(CA[11]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3861 ), .SD(\CODEIF/n3852 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_xnor2x0 \LDCHK/U102  ( .ZN(\LDCHK/n3279 ), .A(\pgmuxout[30] ), .B(
        \pgmuxout[31] ) );
    snl_muxi21x1 \LDIS/U171  ( .ZN(\LDIS/ldexcl[1] ), .A(\LDIS/n3149 ), .B(
        \LDIS/n3150 ), .S(\LDIS/n3134 ) );
    snl_invx1 \PDOSEL/U15  ( .ZN(\PDOSEL/n76 ), .A(SWIT_wire) );
    snl_oai122x0 \LBUS/U581  ( .ZN(ph_timsth), .A(ph_timouth), .B(\LBUS/n1443 
        ), .C(\LBUS/MMBSEL ), .D(LDS), .E(\LBUS/n1442 ) );
    snl_nand13x1 \BLU/U360  ( .ZN(\BLU/n1532 ), .A(\BLU/n1544 ), .B(
        \BLU/n1465 ), .C(\BLU/n1571 ) );
    snl_xor2x0 \CODEIF/U317  ( .Z(\CODEIF/n3960 ), .A(\CODEIF/n3989 ), .B(
        \CODEIF/n3993 ) );
    snl_aoi022x1 \ALUIS/U127  ( .ZN(\ALUIS/n3724 ), .A(\stream4[17] ), .B(
        immbsel), .C(\pk_adb_h[17] ), .D(po_brsel_h) );
    snl_xor2x0 \CODEIF/U330  ( .Z(\CODEIF/n4011 ), .A(CDOUT[17]), .B(CDOUT[22]
        ) );
    snl_aoi012x1 \ALUIS/U100  ( .ZN(\ALUIS/n3749 ), .A(\pgldi[29] ), .B(
        srcbsel), .C(allfbsel) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[4]  ( .Q(\REG_2/RETCNT[4] ), .D(
        \REG_2/ph_retcnt_h[4] ), .EN(\REG_2/n517 ), .RN(\REG_2/n436 ), .SD(
        \REG_2/ncnt2[1] ), .SE(ph_d53lth), .CP(SCLK) );
    snl_nand02x1 \ALUIS/U69  ( .ZN(\pgaluinb[21] ), .A(\ALUIS/n3732 ), .B(
        \ALUIS/n3733 ) );
    snl_invx05 \LDIS/U156  ( .ZN(\LDIS/n3118 ), .A(\pgld32[18] ) );
    snl_mux21x1 \ALUSHT/U25  ( .Z(\pkdptout[26] ), .A(\ALUSHT/pkshtout[26] ), 
        .B(\ALUSHT/pkaluout[26] ), .S(\ALUSHT/n3112 ) );
    snl_invx05 \LBUS/U696  ( .ZN(\LBUS/n1396 ), .A(\LBUS/n1590 ) );
    snl_xor2x0 \CONS/U64  ( .Z(\CONS/n581 ), .A(\CONS/SACO[6] ), .B(
        \pgsdprlh[10] ) );
    snl_nor02x1 \BLU/U347  ( .ZN(\BLU/n1562 ), .A(\BLU/n1559 ), .B(
        \pgbitnoh[2] ) );
    snl_oai012x1 \PDOSEL/U32  ( .ZN(PDH[48]), .A(\PDOSEL/n102 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_and02x1 \SAEXE/U101  ( .Z(\SAEXE/srcread ), .A(\SAEXE/n411 ), .B(
        \SAEXE/singlen ) );
    snl_nand02x1 \PDOSEL/U141  ( .ZN(\PDOSEL/n128 ), .A(CDIN[3]), .B(
        \PDOSEL/n119 ) );
    snl_nor04x0 \LDCHK/U86  ( .ZN(\LDCHK/n3244 ), .A(\LDCHK/n3309 ), .B(
        \pgld32[18] ), .C(\pgld32[5] ), .D(\pgld32[1] ) );
    snl_invx05 \REGF/U812  ( .ZN(\REGF/n8116 ), .A(\pkdptout[11] ) );
    snl_invx05 \REGF/U777  ( .ZN(\REGF/n8186 ), .A(\pgsdprlh[11] ) );
    snl_invx05 \ADOSEL/U70  ( .ZN(\ADOSEL/n4128 ), .A(\pkdptout[29] ) );
    snl_xor2x0 \CODEIF/U245  ( .Z(CPOUT[3]), .A(\CODEIF/n3936 ), .B(
        \CODEIF/n3937 ) );
    snl_xnor2x0 \CONS/U234  ( .ZN(\CONS/n716 ), .A(\pk_idcy_h[22] ), .B(
        \pk_indy_h[22] ) );
    snl_invx05 \BLU/U423  ( .ZN(\BLU/n1530 ), .A(\BLU/n1483 ) );
    snl_oai222x0 \REGF/U485  ( .ZN(\REGF/RI_DPR[8] ), .A(\REGF/n8191 ), .B(
        \REGF/n8160 ), .C(\REGF/n8192 ), .D(\REGF/n8162 ), .E(\REGF/n8126 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U515  ( .Z(\REGF/RI_PCOL[10] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[10]), .C(\stream4[10] ), .D(\REGF/n8209 ) );
    snl_ao2222x1 \REGF/U532  ( .Z(\REGF/RI_SRDA[25] ), .A(PDLIN[25]), .B(
        \ph_pdis_h[9] ), .C(\pgldi[25] ), .D(\REGF/n8210 ), .E(\stream3[25] ), 
        .F(\REGF/n8211 ), .G(\pkdptout[25] ), .H(\REGF/n8212 ) );
    snl_invx05 \REGF/U689  ( .ZN(\REGF/n8084 ), .A(PDLIN[22]) );
    snl_invx05 \REGF/U719  ( .ZN(\REGF/n8133 ), .A(\pgldi[5] ) );
    snl_nor03x0 \LBUS/U673  ( .ZN(\LBUS/n1402 ), .A(\LBUS/n1417 ), .B(
        \LBUS/n1443 ), .C(\LBUS/n1415 ) );
    snl_xor2x0 \CONS/U81  ( .Z(\CONS/n599 ), .A(\pk_pcs1_h[1] ), .B(
        \pk_pc_h[1] ) );
    snl_xor2x0 \CONS/U104  ( .Z(\CONS/n622 ), .A(\pk_idcx_h[7] ), .B(
        \pk_indx_h[7] ) );
    snl_nor02x1 \PDOSEL/U108  ( .ZN(\PDOSEL/n181 ), .A(\pk_pdo_h[8] ), .B(
        \ph_cpudout[8] ) );
    snl_oai122x0 \ADOSEL/U39  ( .ZN(\pgmuxout[28] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4126 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4125 ), .E(
        \ADOSEL/n4151 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[11]  ( .Q(\CODEIF/pfctr[11] ), .D(
        \CODEIF/pfctr415[11] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_muxi21x1 \LDIS/U194  ( .ZN(\LDIS/ldexch[16] ), .A(\LDIS/n3164 ), .B(
        \LDIS/n3163 ), .S(\LDIS/n3165 ) );
    snl_nor03x0 \CONS/U123  ( .ZN(\CONS/n648 ), .A(\CONS/n570 ), .B(
        \CONS/n568 ), .C(\CONS/n569 ) );
    snl_invx05 \CODEIF/U262  ( .ZN(\CODEIF/n3881 ), .A(\CODEIF/pfctr[5] ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[2]  ( .Q(\CODEIF/pfctr[2] ), .D(
        \CODEIF/pfctr415[2] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nor02x1 \LBUS/U654  ( .ZN(\LBUS/n1426 ), .A(\LBUS/n1434 ), .B(
        \LBUS/n1427 ) );
    snl_nand02x1 \BLU/U385  ( .ZN(\BLU/n1507 ), .A(\BLU/n1570 ), .B(
        \BLU/n1568 ) );
    snl_nand13x1 \LBUS/U564  ( .ZN(LDL0), .A(ph_locken_h), .B(\LBUS/n1404 ), 
        .C(\LBUS/ilt[2] ) );
    snl_xnor2x0 \CONS/U213  ( .ZN(\CONS/n695 ), .A(\pk_pc_h[17] ), .B(
        \pk_pcs1_h[17] ) );
    snl_aoi012x1 \BLU/U404  ( .ZN(\BLU/n1575 ), .A(\poalufnc[0] ), .B(
        \BLU/n1519 ), .C(\BLU/n1524 ) );
    snl_and02x1 \REG_2/U142  ( .Z(\ph_cpudout[12] ), .A(\ph_segset_h[12] ), 
        .B(seg_cnfg_h) );
    snl_oai022x1 \REGF/U602  ( .ZN(\REGF/RI_SPR[27] ), .A(\REGF/n8058 ), .B(
        \REGF/n8218 ), .C(\REGF/n8219 ), .D(\REGF/n8153 ) );
    snl_invx05 \REGF/U792  ( .ZN(\REGF/n8143 ), .A(\pkdptout[2] ) );
    snl_invx05 \LDIS/U208  ( .ZN(\LDIS/n3140 ), .A(LIN[22]) );
    snl_nor02x1 \BLU/U329  ( .ZN(\BLU/n1505 ), .A(\BLU/n1541 ), .B(\BLU/n1542 
        ) );
    snl_oai222x0 \REGF/U625  ( .ZN(\REGF/RI_SPR[4] ), .A(\REGF/n8199 ), .B(
        \REGF/n8220 ), .C(\REGF/n8200 ), .D(\REGF/n8221 ), .E(\REGF/n8138 ), 
        .F(\REGF/n8218 ) );
    snl_nand02x1 \ADOSEL/U95  ( .ZN(\ADOSEL/n4148 ), .A(\pgbluext[9] ), .B(
        \ADOSEL/n4156 ) );
    snl_xor2x0 \LDCHK/U44  ( .Z(\LDCHK/n3235 ), .A(\LDCHK/n3256 ), .B(
        \LDCHK/n3257 ) );
    snl_invx05 \CMPX/U29  ( .ZN(\CMPX/n1048 ), .A(ph_lblockh) );
    snl_invx05 \MAIN/U151  ( .ZN(\MAIN/n3632 ), .A(pkaccovf) );
    snl_oai012x1 \LDIS/U138  ( .ZN(\pgldi[24] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3124 ), .C(\LDIS/n3115 ) );
    snl_xor2x0 \LDCHK/U63  ( .Z(\LDCHK/n3263 ), .A(\LDCHK/n3292 ), .B(
        \LDCHK/n3293 ) );
    snl_oai222x0 \REGF/U596  ( .ZN(\REGF/RI_ACC[5] ), .A(\REGF/n8133 ), .B(
        \REGF/n8215 ), .C(\REGF/n8134 ), .D(\REGF/n8216 ), .E(\REGF/n8135 ), 
        .F(\REGF/n8217 ) );
    snl_xnor2x0 \CODEIF/U379  ( .ZN(\CODEIF/n3973 ), .A(CDIN[40]), .B(CDIN[41]
        ) );
    snl_nand02x1 \ALUIS/U149  ( .ZN(\ALUIS/n3662 ), .A(\pk_ada_h[4] ), .B(
        po_arsel_h) );
    snl_invx1 \ALUIS/U20  ( .ZN(\pgaluina[5] ), .A(\ALUIS/n3651 ) );
    snl_ao022x1 \REGF/U421  ( .Z(\REGF/RI_PCOH[12] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[12]), .C(\stream4[44] ), .D(\REGF/n8053 ) );
    snl_invx05 \REGF/U681  ( .ZN(\REGF/n8155 ), .A(PDLIN[29]) );
    snl_invx05 \REGF/U711  ( .ZN(\REGF/n8150 ), .A(PDLIN[0]) );
    snl_invx05 \REGF/U736  ( .ZN(\REGF/n8078 ), .A(PDLIN[24]) );
    snl_oai122x0 \ADOSEL/U31  ( .ZN(\pgmuxout[20] ), .A(\ADOSEL/n4102 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4101 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4143 ) );
    snl_nor02x1 \PDOSEL/U127  ( .ZN(\PDOSEL/n151 ), .A(\pk_pdo_h[16] ), .B(
        \ph_cpudout[16] ) );
    snl_oai122x0 \ADOSEL/U16  ( .ZN(\pgmuxout[5] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4104 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4105 ), .E(
        \ADOSEL/n4106 ) );
    snl_invx05 \PDOSEL/U100  ( .ZN(\PDOSEL/n100 ), .A(CDIN[46]) );
    snl_xor2x0 \CONS/U89  ( .Z(\CONS/n607 ), .A(\pk_idcz_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_aoi012x1 \ALUIS/U84  ( .ZN(\ALUIS/n3705 ), .A(\pgldi[7] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_oai2222x0 \REGF/U362  ( .ZN(\REGF/RI_SRA12M[9] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8123 ), .C(\REGF/n8121 ), .D(\REGF/n8051 ), .E(\REGF/n8189 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8190 ), .H(\REGF/n8230 ) );
    snl_ao2222x1 \REGF/U554  ( .Z(\REGF/RI_SRDA[3] ), .A(PDLIN[3]), .B(
        \ph_pdis_h[9] ), .C(\pgldi[3] ), .D(\REGF/n8210 ), .E(\stream3[3] ), 
        .F(\REGF/n8211 ), .G(\pkdptout[3] ), .H(\REGF/n8212 ) );
    snl_invx05 \REGF/U664  ( .ZN(\REGF/n8185 ), .A(\pgregadrh[11] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[7]  ( .Q(\REGF/RO_LLPSAS[9] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[7] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_xnor2x0 \CODEIF/U371  ( .ZN(\CODEIF/n3964 ), .A(CDIN[54]), .B(CDIN[57]
        ) );
    snl_invx1 \ALUIS/U28  ( .ZN(\pgaluina[7] ), .A(\ALUIS/n3655 ) );
    snl_aoi022x1 \ALUIS/U141  ( .ZN(\ALUIS/n3710 ), .A(\stream4[10] ), .B(
        immbsel), .C(\pk_adb_h[10] ), .D(po_brsel_h) );
    snl_oai022x1 \BLU/U306  ( .ZN(\pkbludgh[10] ), .A(\BLU/n1464 ), .B(
        \BLU/n1480 ), .C(\BLU/n1481 ), .D(\BLU/n1482 ) );
    snl_nand02x1 \CODEIF/U356  ( .ZN(\CODEIF/n3898 ), .A(\CODEIF/pgctrinc[10] 
        ), .B(\CODEIF/n3945 ) );
    snl_ao022x1 \BLUOS/U16  ( .Z(\pgbluext[28] ), .A(\pkbludgh[12] ), .B(
        ph_bit_h), .C(\pkdptout[12] ), .D(ph_word16_h) );
    snl_ao022x1 \LDIS/U117  ( .Z(\pgld16[9] ), .A(\pgld32[9] ), .B(ph_selldl), 
        .C(\pgld32[25] ), .D(ph_selldh) );
    snl_nand02x1 \LDIS/U227  ( .ZN(\LDIS/n3115 ), .A(ph_word16_h), .B(
        \pgld16[15] ) );
    snl_invx05 \SAEXE/U140  ( .ZN(\SAEXE/srcwrit ), .A(\SAEXE/n431 ) );
    snl_ffqrnx1 \LBUS/ilt_reg[4]  ( .Q(\LBUS/ilt[4] ), .D(\LBUS/nlt[4] ), .RN(
        n10734), .CP(SCLK) );
    snl_oai112x0 \PDOSEL/U73  ( .ZN(PDLOUT[0]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n74 ), .C(\PDOSEL/n178 ), .D(\PDOSEL/n179 ) );
    snl_invx05 \MAIN/U159  ( .ZN(\MAIN/n3613 ), .A(\pk_rwrit_h[60] ) );
    snl_oai012x1 \LDIS/U130  ( .ZN(\pgldi[16] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3116 ), .C(\LDIS/n3115 ) );
    snl_mux21x1 \ALUSHT/U43  ( .Z(\pkdptout[0] ), .A(\ALUSHT/pkshtout[0] ), 
        .B(\ALUSHT/pkaluout[0] ), .S(\ALUSHT/n3112 ) );
    snl_ao022x1 \CMPX/U21  ( .Z(ph_word32_h), .A(ph_word32h), .B(ph_saexe_sth), 
        .C(srctype2), .D(\CMPX/n1047 ) );
    snl_xnor2x0 \CONS/U187  ( .ZN(\CONS/n670 ), .A(\pgsdprlh[13] ), .B(
        \CONS/SACO[9] ) );
    snl_oai112x0 \PDOSEL/U54  ( .ZN(PDLOUT[4]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n80 ), .C(\PDOSEL/n132 ), .D(\PDOSEL/n133 ) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[0]  ( .Q(\REG_2/ph_retcnt_h[0] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[0]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_aoi012x1 \BLU/U321  ( .ZN(\BLU/n1517 ), .A(\BLU/n1526 ), .B(
        \BLU/n1527 ), .C(srcbsel) );
    snl_nand02x1 \ALUIS/U166  ( .ZN(\ALUIS/n3676 ), .A(\pk_ada_h[18] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U200  ( .ZN(\LDIS/n3148 ), .A(LIN[18]) );
    snl_ao222x1 \CODEIF/U198  ( .Z(\CODEIF/n3845 ), .A(PA[7]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[4] ), .E(cif_byte), .F(PDLIN[4])
         );
    snl_ao022x1 \MAIN/U137  ( .Z(ph_ebaccwt_h), .A(st_exectl), .B(ph_shelter_h
        ), .C(ebaccsel), .D(ph_filewr_h) );
    snl_aoi112x0 \SAEXE/U109  ( .ZN(ph_dprsel2_h), .A(\SAEXE/n420 ), .B(
        \SAEXE/n421 ), .C(\SAEXE/n422 ), .D(\SAEXE/n423 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[18]  ( .Q(\ph_segset_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[18]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_nand02x1 \ADOSEL/U107  ( .ZN(\ADOSEL/n4133 ), .A(\pgbluext[30] ), .B(
        \ADOSEL/n4156 ) );
    snl_xor2x0 \CODEIF/U338  ( .Z(\CODEIF/n4021 ), .A(CDOUT[3]), .B(CDOUT[1])
         );
    snl_nand02x1 \ALUIS/U61  ( .ZN(\pgaluinb[13] ), .A(\ALUIS/n3716 ), .B(
        \ALUIS/n3717 ) );
    snl_aoi012x1 \ALUIS/U108  ( .ZN(\ALUIS/n3741 ), .A(\pgldi[25] ), .B(
        srcbsel), .C(allfbsel) );
    snl_oai022x1 \REGF/U468  ( .ZN(\REGF/RI_DPR[25] ), .A(\REGF/n8155 ), .B(
        \REGF/n8151 ), .C(\REGF/n8152 ), .D(\REGF/n8156 ) );
    snl_oai222x0 \REGF/U573  ( .ZN(\REGF/RI_ACC[28] ), .A(\REGF/n8065 ), .B(
        \REGF/n8215 ), .C(\REGF/n8066 ), .D(\REGF/n8216 ), .E(\REGF/n8157 ), 
        .F(\REGF/n8217 ) );
    snl_oai022x1 \REGF/U643  ( .ZN(\REGF/RI_TBAI[14] ), .A(\REGF/n8225 ), .B(
        \REGF/n8096 ), .C(\REGF/n8226 ), .D(\REGF/n8171 ) );
    snl_nand02x1 \ALUIS/U46  ( .ZN(\pgaluina[30] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3688 ) );
    snl_and02x1 \UPIF/U14  ( .Z(\ph_pdis_h[8] ), .A(\pk_rread_h[43] ), .B(
        \UPIF/n1046 ) );
    snl_invx05 \LBUS/U589  ( .ZN(LRQ), .A(\LBUS/ilt[0] ) );
    snl_nand13x1 \BLU/U368  ( .ZN(\BLU/n1534 ), .A(\BLU/n1539 ), .B(
        \BLU/n1501 ), .C(\BLU/n1572 ) );
    snl_invx05 \ADOSEL/U78  ( .ZN(\ADOSEL/n4093 ), .A(\pkdptout[1] ) );
    snl_muxi21x1 \LDIS/U179  ( .ZN(\LDIS/ldexch[31] ), .A(\LDIS/n3152 ), .B(
        \LDIS/n3151 ), .S(\LDIS/n3165 ) );
    snl_ao222x1 \CODEIF/U204  ( .Z(\CODEIF/n3851 ), .A(PA[13]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[10] ), .E(cif_byte), .F(PDLIN[10]
        ) );
    snl_oai122x0 \CODEIF/U223  ( .ZN(\CODEIF/pfctr415[2] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3872 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3873 ), .E(
        \CODEIF/n3874 ) );
    snl_oa022x1 \LBUS/U615  ( .Z(\LBUS/n1398 ), .A(\LBUS/n1461 ), .B(
        \LBUS/n1462 ), .C(\LBUS/n1453 ), .D(\LBUS/n1591 ) );
    snl_nor04x0 \CONS/U162  ( .ZN(\CONS/n344 ), .A(\CONS/n746 ), .B(
        \CONS/n636 ), .C(\CONS/n634 ), .D(\CONS/n635 ) );
    snl_xnor2x0 \CONS/U252  ( .ZN(\CONS/n736 ), .A(\pk_idcx_h[21] ), .B(
        \pk_indx_h[21] ) );
    snl_nand13x1 \BLU/U445  ( .ZN(\BLU/n1585 ), .A(po_cmfsel_h), .B(
        \BLU/n1558 ), .C(pkaluopc) );
    snl_xnor2x0 \CONS/U275  ( .ZN(\CONS/n340 ), .A(\pk_idcw_h[5] ), .B(
        \pk_indw_h[5] ) );
    snl_xnor2x0 \CODEIF/U394  ( .ZN(\CODEIF/n3988 ), .A(CDIN[9]), .B(CDIN[12])
         );
    snl_xnor2x0 \CODEIF/U415  ( .ZN(\CODEIF/n4041 ), .A(CDOUT[26]), .B(CDOUT
        [27]) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[22]  ( .Q(\pgld32[22] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[22] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_oai222x0 \REGF/U473  ( .ZN(\REGF/RI_DPR[20] ), .A(\REGF/n8167 ), .B(
        \REGF/n8160 ), .C(\REGF/n8168 ), .D(\REGF/n8162 ), .E(\REGF/n8090 ), 
        .F(\REGF/n8151 ) );
    snl_invx05 \REGF/U743  ( .ZN(\REGF/n8094 ), .A(\pgldi[18] ) );
    snl_invx05 \REGF/U758  ( .ZN(\REGF/n8200 ), .A(\pgsdprlh[4] ) );
    snl_sffqenrnx1 \MAIN/accovf_reg  ( .Q(\MAIN/accovf ), .D(1'b0), .EN(1'b1), 
        .RN(\MAIN/n3611 ), .SD(\MAIN/*cell*4603/U7/CONTROL1 ), .SE(
        \MAIN/*cell*4603/U16/CONTROL1 ), .CP(SCLK) );
    snl_and08x1 \CONS/U145  ( .Z(\CONS/n535 ), .A(\CONS/n703 ), .B(\CONS/n704 
        ), .C(\CONS/n705 ), .D(\CONS/n706 ), .E(\CONS/n707 ), .F(\CONS/n708 ), 
        .G(\CONS/n709 ), .H(\CONS/n702 ) );
    snl_invx05 \PDOSEL/U96  ( .ZN(\PDOSEL/n104 ), .A(CDIN[50]) );
    snl_nand02x1 \PDOSEL/U149  ( .ZN(\PDOSEL/n158 ), .A(CDIN[21]), .B(
        \PDOSEL/n119 ) );
    snl_nor02x1 \LBUS/U629  ( .ZN(\LBUS/n1597 ), .A(pgldperrh), .B(LBER) );
    snl_oa012x1 \LBUS/U632  ( .Z(\LBUS/n1446 ), .A(\LBUS/n1409 ), .B(
        \LBUS/n1445 ), .C(\LBUS/n1431 ) );
    snl_nand12x1 \ADOSEL/U44  ( .ZN(\ADOSEL/n4087 ), .A(\ADOSEL/n4155 ), .B(
        ph_word32_h) );
    snl_bufx1 \ALUIS/U6  ( .Z(\pgaluina[3] ), .A(\ALUIS/n3754 ) );
    snl_oai012x1 \LDCHK/U95  ( .ZN(\LDCHK/n3236 ), .A(\LDCHK/n3253 ), .B(
        \LDCHK/n3268 ), .C(ph_pdhen_h) );
    snl_nand02x1 \PDOSEL/U152  ( .ZN(\PDOSEL/n120 ), .A(CDIN[1]), .B(
        \PDOSEL/n119 ) );
    snl_invx1 \LDIS/U97  ( .ZN(\LDIS/n3113 ), .A(ph_word32_h) );
    snl_invx05 \REGF/U801  ( .ZN(\REGF/n8086 ), .A(\pkdptout[21] ) );
    snl_oai2222x0 \REGF/U379  ( .ZN(\REGF/RI_SRA12M[13] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8111 ), .C(\REGF/n8109 ), .D(\REGF/n8051 ), .E(\REGF/n8181 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8182 ) );
    snl_oai222x0 \REGF/U454  ( .ZN(\REGF/RI_EACC[11] ), .A(\REGF/n8115 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8116 ), .E(\REGF/n8117 ), 
        .F(\REGF/n8059 ) );
    snl_or08x1 \REGF/U658  ( .Z(\REGF/RO_PSTA[16] ), .A(\REGF/RO_EST1[3] ), 
        .B(\REGF/RO_EST1[1] ), .C(\REGF/RO_EST1[7] ), .D(\REGF/RO_EST1[2] ), 
        .E(\REGF/RO_EST1[5] ), .F(\REGF/RO_EST1[6] ), .G(\REGF/RO_EST1[0] ), 
        .H(\REGF/RO_EST1[4] ) );
    snl_invx05 \REGF/U764  ( .ZN(\REGF/n8164 ), .A(\pgsdprlh[22] ) );
    snl_aoi022x1 \REGF/U826  ( .ZN(\REGF/n8214 ), .A(\pkdptout[0] ), .B(
        \REGF/n8212 ), .C(\stream3[0] ), .D(\REGF/n8211 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[11]  ( .Q(\ph_segset_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[11]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_oai122x0 \CODEIF/U238  ( .ZN(\CODEIF/pfctr415[17] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3917 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3918 ), .E(
        \CODEIF/n3919 ) );
    snl_mux21x1 \SHTCD/U15  ( .Z(\phshtd[1] ), .A(\pgld16[1] ), .B(
        \stream4[1] ), .S(immbsel) );
    snl_xnor2x0 \CONS/U249  ( .ZN(\CONS/n728 ), .A(\pk_idcx_h[8] ), .B(
        \pk_indx_h[8] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[22]  ( .Q(\ph_segset_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[22]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[10]  ( .Q(\REGF/RO_LLPSAS[14] ), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[10] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_nand02x1 \ADOSEL/U63  ( .ZN(\ADOSEL/n4138 ), .A(ph_word32_h), .B(
        \ADOSEL/n4157 ) );
    snl_xnor2x0 \CONS/U179  ( .ZN(\CONS/n662 ), .A(\pgsdprlh[18] ), .B(
        \pk_saco_lh[18] ) );
    snl_invx05 \LDIS/U162  ( .ZN(\LDIS/n3116 ), .A(\pgld32[16] ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[15]  ( .Q(\pgld32[15] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexcl[15] ), .SE(lo_data_lth), .CP(SCLK
        ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[18]  ( .Q(\pgld32[18] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[18] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_xor2x0 \CODEIF/U294  ( .Z(\CODEIF/n3924 ), .A(\CODEIF/n3955 ), .B(
        \CODEIF/n3956 ) );
    snl_or02x1 \ALUSHT/U11  ( .Z(pkaluovf), .A(\ALUSHT/slaovf ), .B(
        \ALUSHT/aluovf ) );
    snl_xor2x0 \CONS/U50  ( .Z(\CONS/n572 ), .A(\pgsdprlh[23] ), .B(
        \pk_saco_lh[23] ) );
    snl_nand03x0 \SAEXE/U135  ( .ZN(\SAEXE/n421 ), .A(ph_saexe_sth), .B(
        \SAEXE/n411 ), .C(\SAEXE/sequen ) );
    snl_xor2x0 \CODEIF/U304  ( .Z(\CODEIF/n3971 ), .A(CDIN[45]), .B(CDIN[46])
         );
    snl_nand02x1 \BLU/U373  ( .ZN(\BLU/n1492 ), .A(\BLU/n1569 ), .B(
        \BLU/n1561 ) );
    snl_aoi012x1 \ALUIS/U134  ( .ZN(\ALUIS/n3717 ), .A(\pgldi[13] ), .B(
        srcbsel), .C(allfbsel) );
    snl_xnor2x0 \LDCHK/U111  ( .ZN(\LDCHK/n3288 ), .A(\pgmuxout[14] ), .B(
        \pgmuxout[15] ) );
    snl_and02x1 \LBUS/U592  ( .Z(ph_srdalth), .A(\LBUS/srdalth ), .B(
        \LBUS/n1404 ) );
    snl_and02x1 \REGF/U568  ( .Z(\REGF/RO_LPSAS2156[10] ), .A(ph_tirtendh), 
        .B(ph_sastlth) );
    snl_xor2x0 \CODEIF/U323  ( .Z(\CODEIF/n4000 ), .A(CDOUT[48]), .B(CDOUT[46]
        ) );
    snl_aoi022x1 \ALUIS/U113  ( .ZN(\ALUIS/n3736 ), .A(\stream4[23] ), .B(
        immbsel), .C(\pk_adb_h[23] ), .D(po_brsel_h) );
    snl_ffandx1 \MAIN/EXCEP_1H_reg  ( .Q(\MAIN/EXCEP_1H ), .A(pk_excp_h), .B(
        \MAIN/sw_end ), .CP(SCLK) );
    snl_nor02x1 \BLU/U354  ( .ZN(\BLU/n1569 ), .A(\BLU/n1566 ), .B(
        \pgbitnoh[3] ) );
    snl_ao022x1 \REGF/U428  ( .Z(\REGF/RI_PCOH[5] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[5]), .C(\stream4[37] ), .D(\REGF/n8053 ) );
    snl_ao022x1 \REGF/U496  ( .Z(\REGF/RI_PCOL[29] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[29]), .C(\stream4[29] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U506  ( .Z(\REGF/RI_PCOL[19] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[19]), .C(\stream4[19] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U521  ( .Z(\REGF/RI_PCOL[4] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[4]), .C(\stream4[4] ), .D(\REGF/n8209 ) );
    snl_and02x1 \ALUIS/U14  ( .Z(\ALUIS/n3647 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3669 ) );
    snl_xor2x0 \LDCHK/U39  ( .Z(\LDCHK/n3250 ), .A(\LDCHK/n3251 ), .B(
        \LDCHK/n3252 ) );
    snl_oai012x1 \LDIS/U145  ( .ZN(\pgldi[31] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3131 ), .C(\LDIS/n3115 ) );
    snl_oai012x1 \PDOSEL/U21  ( .ZN(PDH[37]), .A(\PDOSEL/n81 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_or03x1 \SAEXE/U112  ( .Z(phrelbsth), .A(\SAEXE/sa_start1 ), .B(
        \SAEXE/sa_start2 ), .C(\SAEXE/sa_start3 ) );
    snl_mux21x1 \ALUSHT/U36  ( .Z(\pkdptout[16] ), .A(\ALUSHT/pkshtout[16] ), 
        .B(\ALUSHT/pkaluout[16] ), .S(\ALUSHT/n3112 ) );
    snl_and02x1 \LBUS/U685  ( .Z(\LBUS/n1412 ), .A(\LBUS/n1611 ), .B(
        \LBUS/n1608 ) );
    snl_xor2x0 \CONS/U77  ( .Z(\CONS/n595 ), .A(\pk_pcs1_h[16] ), .B(
        \pk_pc_h[16] ) );
    snl_oai222x0 \REGF/U611  ( .ZN(\REGF/RI_SPR[18] ), .A(\REGF/n8171 ), .B(
        \REGF/n8220 ), .C(\REGF/n8172 ), .D(\REGF/n8221 ), .E(\REGF/n8096 ), 
        .F(\REGF/n8218 ) );
    snl_and12x1 \REGF/U781  ( .Z(\REGF/n8209 ), .A(\ph_pdis_h[6] ), .B(
        ph_rgfile_h) );
    snl_nand02x1 \ADOSEL/U86  ( .ZN(\ADOSEL/n4103 ), .A(\pgbluext[4] ), .B(
        \ADOSEL/n4156 ) );
    snl_or02x1 \MAIN/U142  ( .Z(\MAIN/dprw_inhibith ), .A(\MAIN/dprw_tap2 ), 
        .B(\MAIN/dprw_tap1 ) );
    snl_xor2x0 \LDCHK/U57  ( .Z(\LDCHK/n3257 ), .A(\LDCHK/n3280 ), .B(
        \LDCHK/n3281 ) );
    snl_oai022x1 \REGF/U636  ( .ZN(\REGF/RI_TBAI[23] ), .A(\REGF/n8225 ), .B(
        \REGF/n8058 ), .C(\REGF/n8226 ), .D(\REGF/n8153 ) );
    snl_invx05 \MAIN/U165  ( .ZN(\MAIN/n3619 ), .A(ph_exstgb_h) );
    snl_oai112x0 \PDOSEL/U68  ( .ZN(PDLOUT[21]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n107 ), .C(\PDOSEL/n158 ), .D(\PDOSEL/n159 ) );
    snl_nand02x1 \ALUIS/U33  ( .ZN(\pgaluina[17] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3675 ) );
    snl_xor2x0 \LDCHK/U70  ( .Z(\LDCHK/n3252 ), .A(\LDCHK/n3298 ), .B(
        \LDCHK/n3299 ) );
    snl_invx05 \CODEIF/U256  ( .ZN(\CODEIF/n3890 ), .A(\CODEIF/pfctr[8] ) );
    snl_ffqsnx1 \LBUS/l_pd_reg  ( .Q(LPDOUT), .D(
        \LBUS/*cell*3982/U111/CONTROL2 ), .SN(n10734), .CP(SCLK) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[5]  ( .Q(\pgld32[5] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[5] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_invx05 \LBUS/U660  ( .ZN(\LBUS/*cell*3982/U70/CONTROL1 ), .A(
        \LBUS/n1414 ) );
    snl_xnor2x0 \CONS/U227  ( .ZN(\CONS/n533 ), .A(\pk_idcz_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_nand04x0 \BLU/U430  ( .ZN(\BLU/n1518 ), .A(pk_bitdatah), .B(
        \BLU/n1527 ), .C(srcbsel), .D(\BLU/n1586 ) );
    snl_nand02x1 \LBUS/U647  ( .ZN(\LBUS/n1430 ), .A(\LBUS/ilt[2] ), .B(
        \LBUS/n1452 ) );
    snl_xor2x0 \CONS/U92  ( .Z(\CONS/n610 ), .A(\pk_idcy_h[3] ), .B(
        \pk_indy_h[3] ) );
    snl_xor2x0 \CONS/U117  ( .Z(\CONS/n635 ), .A(\pk_idcw_h[7] ), .B(
        \pk_indw_h[7] ) );
    snl_invx05 \CODEIF/U271  ( .ZN(\CODEIF/n3870 ), .A(PDLIN[1]) );
    snl_muxi21x1 \LDIS/U187  ( .ZN(\LDIS/ldexch[23] ), .A(\LDIS/n3138 ), .B(
        \LDIS/n3137 ), .S(\LDIS/n3165 ) );
    snl_and02x1 \LBUS/U577  ( .Z(ph_lbaovf), .A(\LBUS/n1435 ), .B(\LBUS/n1436 
        ) );
    snl_nand04x0 \CONS/U130  ( .ZN(\CONS/n566 ), .A(\CONS/n668 ), .B(
        \CONS/n669 ), .C(\CONS/n667 ), .D(\CONS/n670 ) );
    snl_and02x1 \REG_2/U151  ( .Z(\ph_cpudout[21] ), .A(\ph_segset_h[21] ), 
        .B(seg_cnfg_h) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[26]  ( .Q(\pgld32[26] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[26] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_xnor2x0 \CONS/U200  ( .ZN(\CONS/n684 ), .A(\pk_pc_h[18] ), .B(
        \pk_pcs2_h[18] ) );
    snl_invx05 \BLU/U396  ( .ZN(\BLU/n1479 ), .A(\pgld16[11] ) );
    snl_invx05 \BLU/U417  ( .ZN(\BLU/n1541 ), .A(\BLU/n1507 ) );
    snl_invx05 \REGF/U688  ( .ZN(\REGF/n8163 ), .A(\pgregadrh[22] ) );
    snl_xor2x0 \CODEIF/U244  ( .Z(\CODEIF/n3933 ), .A(\CODEIF/n3934 ), .B(
        \CODEIF/n3935 ) );
    snl_xnor2x0 \CONS/U235  ( .ZN(\CONS/n715 ), .A(\pk_idcy_h[12] ), .B(
        \pk_indy_h[12] ) );
    snl_invx05 \BLU/U422  ( .ZN(\BLU/n1538 ), .A(\BLU/n1489 ) );
    snl_nand13x1 \LBUS/U672  ( .ZN(\LBUS/n1608 ), .A(\LBUS/word32odphase ), 
        .B(\LBUS/n1457 ), .C(ph_word32_h) );
    snl_xor2x0 \CONS/U80  ( .Z(\CONS/n598 ), .A(\pk_pcs1_h[2] ), .B(
        \pk_pc_h[2] ) );
    snl_invx05 \REGF/U718  ( .ZN(\REGF/n8130 ), .A(\pgldi[6] ) );
    snl_oai222x0 \REGF/U446  ( .ZN(\REGF/RI_EACC[19] ), .A(\REGF/n8091 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8092 ), .E(\REGF/n8093 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U461  ( .ZN(\REGF/RI_EACC[4] ), .A(\REGF/n8136 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8137 ), .E(\REGF/n8138 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U484  ( .ZN(\REGF/RI_DPR[9] ), .A(\REGF/n8189 ), .B(
        \REGF/n8160 ), .C(\REGF/n8190 ), .D(\REGF/n8162 ), .E(\REGF/n8123 ), 
        .F(\REGF/n8151 ) );
    snl_ao2222x1 \REGF/U533  ( .Z(\REGF/RI_SRDA[24] ), .A(PDLIN[24]), .B(
        \ph_pdis_h[9] ), .C(\pgldi[24] ), .D(\REGF/n8210 ), .E(\stream3[24] ), 
        .F(\REGF/n8211 ), .G(\pkdptout[24] ), .H(\REGF/n8212 ) );
    snl_oai122x0 \ADOSEL/U38  ( .ZN(\pgmuxout[27] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4123 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4122 ), .E(
        \ADOSEL/n4150 ) );
    snl_invx05 \LDIS/U195  ( .ZN(\LDIS/n3163 ), .A(LIN[0]) );
    snl_aoi122x0 \LBUS/U655  ( .ZN(\LBUS/n1449 ), .A(\LBUS/n1606 ), .B(
        \LBUS/ilt[2] ), .C(\LBUS/n1607 ), .D(\LBUS/n1452 ), .E(\LBUS/n1598 )
         );
    snl_xor2x0 \CONS/U105  ( .Z(\CONS/n623 ), .A(\pk_idcx_h[1] ), .B(
        \pk_indx_h[1] ) );
    snl_nor02x1 \PDOSEL/U109  ( .ZN(\PDOSEL/n147 ), .A(\pk_pdo_h[7] ), .B(
        \ph_cpudout[7] ) );
    snl_nand02x1 \CONS/U122  ( .ZN(\CONS/n647 ), .A(\CONS/n298 ), .B(
        \CONS/n300 ) );
    snl_invx05 \CODEIF/U263  ( .ZN(\CODEIF/n3882 ), .A(PDLIN[5]) );
    snl_nand02x1 \LBUS/U565  ( .ZN(\LBUS/*cell*3982/U176/CONTROL1 ), .A(
        \LBUS/n1405 ), .B(\LBUS/n1401 ) );
    snl_xnor2x0 \CONS/U212  ( .ZN(\CONS/n696 ), .A(\pk_pc_h[12] ), .B(
        \pk_pcs1_h[12] ) );
    snl_nor02x1 \BLU/U405  ( .ZN(\BLU/n1576 ), .A(\BLU/n1522 ), .B(\BLU/n1523 
        ) );
    snl_invx05 \LDIS/U209  ( .ZN(\LDIS/n3137 ), .A(LIN[7]) );
    snl_and02x1 \REG_2/U143  ( .Z(\ph_cpudout[13] ), .A(\ph_segset_h[13] ), 
        .B(seg_cnfg_h) );
    snl_invx05 \BLU/U384  ( .ZN(\BLU/n1509 ), .A(\pgld16[1] ) );
    snl_nor02x1 \BLU/U328  ( .ZN(\BLU/n1502 ), .A(\BLU/n1539 ), .B(\BLU/n1540 
        ) );
    snl_oai022x1 \REGF/U603  ( .ZN(\REGF/RI_SPR[26] ), .A(\REGF/n8062 ), .B(
        \REGF/n8218 ), .C(\REGF/n8219 ), .D(\REGF/n8154 ) );
    snl_nand02x1 \ADOSEL/U94  ( .ZN(\ADOSEL/n4149 ), .A(\pgbluext[26] ), .B(
        \ADOSEL/n4156 ) );
    snl_ao022x1 \CMPX/U28  ( .Z(ph_atchkenh), .A(phatchkh), .B(ph_saexe_sth), 
        .C(po_atchk_h), .D(\CMPX/n1047 ) );
    snl_invx05 \MAIN/U150  ( .ZN(\MAIN/n3618 ), .A(stage_b) );
    snl_oai012x1 \LDIS/U139  ( .ZN(\pgldi[25] ), .A(\LDIS/n3125 ), .B(
        \LDIS/n3113 ), .C(\LDIS/n3115 ) );
    snl_oai222x0 \REGF/U624  ( .ZN(\REGF/RI_SPR[5] ), .A(\REGF/n8197 ), .B(
        \REGF/n8220 ), .C(\REGF/n8198 ), .D(\REGF/n8221 ), .E(\REGF/n8135 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U793  ( .ZN(\REGF/n8064 ), .A(\pkdptout[29] ) );
    snl_xor2x0 \LDCHK/U45  ( .Z(\LDCHK/n3234 ), .A(\LDCHK/n3258 ), .B(
        \LDCHK/n3259 ) );
    snl_xor2x0 \LDCHK/U62  ( .Z(\LDCHK/n3262 ), .A(\LDCHK/n3290 ), .B(
        \LDCHK/n3291 ) );
    snl_xnor2x0 \CODEIF/U378  ( .ZN(\CODEIF/n3972 ), .A(CDIN[39]), .B(CDIN[42]
        ) );
    snl_nand02x2 \ALUIS/U21  ( .ZN(\pgaluina[8] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3666 ) );
    snl_nand02x1 \ALUIS/U148  ( .ZN(\ALUIS/n3663 ), .A(\pk_ada_h[5] ), .B(
        po_arsel_h) );
    snl_ao022x1 \REGF/U514  ( .Z(\REGF/RI_PCOL[11] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[11]), .C(\stream4[11] ), .D(\REGF/n8209 ) );
    snl_invx05 \REGF/U751  ( .ZN(\REGF/n8118 ), .A(\pgldi[10] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[3]  ( .Q(\REGF/RO_LLPSAS[5] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[3] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_invx05 \CODEIF/U286  ( .ZN(\CODEIF/n3899 ), .A(\CODEIF/pfctr[11] ) );
    snl_xor2x0 \CODEIF/U316  ( .Z(\CODEIF/n3992 ), .A(CDIN[3]), .B(CDIN[5]) );
    snl_invx05 \MAIN/U119  ( .ZN(\MAIN/n3610 ), .A(n10731) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[4]  ( .Q(\REG_2/ph_retcnt_h[4] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[4]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_muxi21x1 \LDIS/U170  ( .ZN(\LDIS/ldexcl[2] ), .A(\LDIS/n3147 ), .B(
        \LDIS/n3148 ), .S(\LDIS/n3134 ) );
    snl_nand03x2 \PDOSEL/U14  ( .ZN(\PDOSEL/n114 ), .A(SWIT_wire), .B(PA02), 
        .C(code_area_h) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[8]  ( .Q(\pgld32[8] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[8] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_nand02x1 \CONS/U42  ( .ZN(\CONS/n549 ), .A(\CONS/n557 ), .B(
        \CONS/n558 ) );
    snl_nor04x0 \SAEXE/U127  ( .ZN(ph_bitsrch), .A(\SAEXE/n413 ), .B(
        \pk_psae_h[0] ), .C(\pk_psae_h[1] ), .D(\pk_psae_h[7] ) );
    snl_aoi012x1 \ALUIS/U126  ( .ZN(\ALUIS/n3725 ), .A(\pgldi[17] ), .B(
        srcbsel), .C(allfbsel) );
    snl_xnor2x0 \LDCHK/U103  ( .ZN(\LDCHK/n3280 ), .A(\pgmuxout[24] ), .B(
        \pgmuxout[25] ) );
    snl_nand13x1 \BLU/U361  ( .ZN(\BLU/n1529 ), .A(\BLU/n1532 ), .B(
        \BLU/n1477 ), .C(\BLU/n1486 ) );
    snl_oai012x1 \LBUS/U580  ( .ZN(ph_initldh), .A(\LBUS/n1395 ), .B(
        \LBUS/n1396 ), .C(\LBUS/n1442 ) );
    snl_xor2x0 \CODEIF/U331  ( .Z(\CODEIF/n4012 ), .A(CDOUT[20]), .B(
        \CODEIF/n4011 ) );
    snl_nor02x1 \BLU/U346  ( .ZN(\BLU/n1561 ), .A(\BLU/n1560 ), .B(
        \pgbitnoh[0] ) );
    snl_nand02x1 \ALUIS/U68  ( .ZN(\pgaluinb[20] ), .A(\ALUIS/n3730 ), .B(
        \ALUIS/n3731 ) );
    snl_aoi022x1 \ALUIS/U101  ( .ZN(\ALUIS/n3748 ), .A(\stream4[29] ), .B(
        immbsel), .C(\pk_adb_h[29] ), .D(po_brsel_h) );
    snl_nor04x0 \LDCHK/U87  ( .ZN(\LDCHK/n3241 ), .A(\pgld32[17] ), .B(
        \pgld32[25] ), .C(\pgld32[3] ), .D(\pgld32[26] ) );
    snl_invx05 \LDIS/U157  ( .ZN(\LDIS/n3129 ), .A(\pgld32[29] ) );
    snl_ffqrnx1 \LBUS/ilt_reg[0]  ( .Q(\LBUS/ilt[0] ), .D(\LBUS/nlt[0] ), .RN(
        n10734), .CP(SCLK) );
    snl_oai012x1 \PDOSEL/U33  ( .ZN(PDH[49]), .A(\PDOSEL/n103 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_mux21x1 \ALUSHT/U24  ( .Z(\pkdptout[27] ), .A(\ALUSHT/pkshtout[27] ), 
        .B(\ALUSHT/pkaluout[27] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U65  ( .Z(\CONS/n582 ), .A(\pgsdprlh[9] ), .B(
        \CONS/SACO[5] ) );
    snl_oa012x1 \SAEXE/U100  ( .Z(\SAEXE/*cell*3651/U4/CONTROL1 ), .A(
        \SAEXE/adovflth2 ), .B(\SAEXE/adovflth1 ), .C(pgadrovfh) );
    snl_invx05 \REGF/U813  ( .ZN(\REGF/n8119 ), .A(\pkdptout[10] ) );
    snl_invx05 \ADOSEL/U56  ( .ZN(\ADOSEL/n4101 ), .A(\pkdptout[20] ) );
    snl_nand02x1 \PDOSEL/U140  ( .ZN(\PDOSEL/n132 ), .A(CDIN[4]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \REGF/U834  ( .ZN(\REGF/n8233 ), .A(po_imdselh) );
    snl_invx05 \REGF/U776  ( .ZN(\REGF/n8184 ), .A(\pgsdprlh[12] ) );
    snl_invx05 \REGF/U808  ( .ZN(\REGF/n8104 ), .A(\pkdptout[15] ) );
    snl_invx05 \ADOSEL/U71  ( .ZN(\ADOSEL/n4126 ), .A(\pkdptout[12] ) );
    snl_nor02x2 \CODEIF/U216  ( .ZN(\CODEIF/n3929 ), .A(cif_byte), .B(cif_cont
        ) );
    snl_oai122x0 \CODEIF/U231  ( .ZN(\CODEIF/pfctr415[10] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3896 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3897 ), .E(
        \CODEIF/n3898 ) );
    snl_invx05 \LBUS/U607  ( .ZN(\LBUS/n1452 ), .A(\LBUS/ilt[4] ) );
    snl_xnor2x0 \CONS/U170  ( .ZN(\CONS/n554 ), .A(\pk_saco_hh[29] ), .B(
        \pgsdprhh[29] ) );
    snl_xnor2x0 \CODEIF/U386  ( .ZN(\CODEIF/n3981 ), .A(CDIN[25]), .B(CDIN[26]
        ) );
    snl_xnor2x0 \CODEIF/U420  ( .ZN(\CODEIF/n4017 ), .A(CDOUT[11]), .B(CDOUT
        [13]) );
    snl_xnor2x0 \CONS/U240  ( .ZN(\CONS/n524 ), .A(\pk_idcy_h[6] ), .B(
        \pk_indy_h[6] ) );
    snl_ao022x1 \REG_2/U136  ( .Z(\ph_cpudout[6] ), .A(\ph_segset_h[6] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[6] ), .D(ret_cont_h) );
    snl_xnor2x0 \CODEIF/U407  ( .ZN(\CODEIF/n4002 ), .A(CDOUT[40]), .B(CDOUT
        [42]) );
    snl_xnor2x0 \CONS/U267  ( .ZN(\CONS/n748 ), .A(\pk_idcw_h[16] ), .B(
        \pk_indw_h[16] ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[1]  ( .Q(\pgld32[1] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[1] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_nor04x0 \CONS/U157  ( .ZN(\CONS/n518 ), .A(\CONS/n734 ), .B(
        \CONS/n627 ), .C(\CONS/n625 ), .D(\CONS/n626 ) );
    snl_invx05 \PDOSEL/U84  ( .ZN(\PDOSEL/n79 ), .A(CDIN[35]) );
    snl_oai2222x0 \REGF/U357  ( .ZN(\REGF/RI_SRA12M[18] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8096 ), .C(\REGF/n8094 ), .D(\REGF/n8051 ), .E(\REGF/n8171 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8172 ) );
    snl_invx05 \REGF/U676  ( .ZN(\REGF/n8153 ), .A(\pgsdprhh[31] ) );
    snl_nor08x1 \LDCHK/U30  ( .ZN(\LDCHK/n3230 ), .A(\pgld32[16] ), .B(
        \pgld32[24] ), .C(\pgld32[8] ), .D(\pgld32[11] ), .E(\pgld32[15] ), 
        .F(\pgld32[14] ), .G(\pgld32[23] ), .H(\pgld32[6] ) );
    snl_invx05 \LBUS/U620  ( .ZN(\LBUS/n1438 ), .A(ph_rmw2h) );
    snl_nor02x1 \MAIN/U125  ( .ZN(\MAIN/n3616 ), .A(ph_cperr_h), .B(
        \MAIN/exe_end ) );
    snl_oai012x1 \PDOSEL/U28  ( .ZN(PDH[44]), .A(\PDOSEL/n98 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_oai022x1 \REGF/U370  ( .ZN(\REGF/RI_TBAI[22] ), .A(\REGF/n8225 ), .B(
        \REGF/n8062 ), .C(\REGF/n8226 ), .D(\REGF/n8154 ) );
    snl_ao2222x1 \REGF/U546  ( .Z(\REGF/RI_SRDA[11] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[11]), .C(\pgldi[11] ), .D(\REGF/n8210 ), .E(\stream3[11] ), .F(
        \REGF/n8211 ), .G(\pkdptout[11] ), .H(\REGF/n8212 ) );
    snl_and02x1 \REGF/U561  ( .Z(\REGF/RO_LPSAS2156[3] ), .A(ph_sastlth), .B(
        \REGF/RO_EST1[5] ) );
    snl_nand02x1 \ALUIS/U73  ( .ZN(\pgaluinb[25] ), .A(\ALUIS/n3740 ), .B(
        \ALUIS/n3741 ) );
    snl_xor2x0 \LDCHK/U118  ( .Z(\LDCHK/n3248 ), .A(\LDCHK/n3297 ), .B(
        \pgld32[3] ) );
    snl_nand02x3 \REGF/U395  ( .ZN(\REGF/n8215 ), .A(po_ldis_h), .B(
        \REGF/n8217 ) );
    snl_ao022x1 \REGF/U414  ( .Z(\REGF/RI_PCOH[19] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[19]), .C(\stream4[51] ), .D(\REGF/n8053 ) );
    snl_ao2222x1 \REGF/U528  ( .Z(\REGF/RI_SRDA[29] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[29]), .C(\pgldi[29] ), .D(\REGF/n8210 ), .E(\stream3[29] ), .F(
        \REGF/n8211 ), .G(\pkdptout[29] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U618  ( .ZN(\REGF/RI_SPR[11] ), .A(\REGF/n8185 ), .B(
        \REGF/n8220 ), .C(\REGF/n8186 ), .D(\REGF/n8221 ), .E(\REGF/n8117 ), 
        .F(\REGF/n8218 ) );
    snl_oai022x1 \REGF/U651  ( .ZN(\REGF/RI_TBAI[3] ), .A(\REGF/n8225 ), .B(
        \REGF/n8129 ), .C(\REGF/n8226 ), .D(\REGF/n8193 ) );
    snl_nand02x1 \ALUIS/U54  ( .ZN(\pgaluinb[6] ), .A(\ALUIS/n3702 ), .B(
        \ALUIS/n3703 ) );
    snl_ffqrnx1 \MAIN/dprw_tap2_reg  ( .Q(\MAIN/dprw_tap2 ), .D(
        \MAIN/dprw_tap1 ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_xor2x0 \CODEIF/U363  ( .Z(\CODEIF/n4024 ), .A(\CODEIF/n4025 ), .B(
        \CODEIF/n4006 ) );
    snl_mux21x1 \ALUSHT/U18  ( .Z(\pkdptout[3] ), .A(\ALUSHT/pkshtout[3] ), 
        .B(\ALUSHT/pkaluout[3] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U59  ( .Z(\CONS/n576 ), .A(\pgsdprlh[6] ), .B(
        \CONS/SACO[2] ) );
    snl_oai022x1 \BLU/U314  ( .ZN(\pkbludgh[2] ), .A(\BLU/n1464 ), .B(
        \BLU/n1504 ), .C(\BLU/n1505 ), .D(\BLU/n1506 ) );
    snl_nand02x1 \ALUIS/U153  ( .ZN(\ALUIS/n3660 ), .A(\pk_ada_h[2] ), .B(
        po_arsel_h) );
    snl_oai023x2 \SAEXE/U98  ( .ZN(ph_srcadr2_h), .A(\SAEXE/n421 ), .B(
        \pk_psae_h[4] ), .C(\SAEXE/n423 ), .D(\SAEXE/n413 ), .E(\SAEXE/n425 )
         );
    snl_ao022x1 \BLUOS/U23  ( .Z(\pgbluext[4] ), .A(\pkbludgh[4] ), .B(
        ph_bit_h), .C(\pkdptout[4] ), .D(ph_word16_h) );
    snl_nor02x1 \CONS/U37  ( .ZN(\CONS/n547 ), .A(ph_wrdsrc_h), .B(ph_bitsrc_h
        ) );
    snl_xor2x0 \LDCHK/U79  ( .Z(\LDCHK/n3306 ), .A(\pgld32[24] ), .B(
        \pgld32[25] ) );
    snl_ao022x1 \LDIS/U105  ( .Z(\pgld16[3] ), .A(ph_selldl), .B(\pgld32[3] ), 
        .C(ph_selldh), .D(\pgld32[19] ) );
    snl_or02x1 \CMPX/U14  ( .Z(ph_bnolt_h), .A(phbnolth), .B(pgbnolth) );
    snl_oai112x0 \PDOSEL/U61  ( .ZN(PDLOUT[7]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n92 ), .C(\PDOSEL/n146 ), .D(\PDOSEL/n147 ) );
    snl_invx05 \REGF/U788  ( .ZN(\REGF/n8137 ), .A(\pkdptout[4] ) );
    snl_ao022x1 \LDIS/U122  ( .Z(\pgldi[12] ), .A(ph_word32_h), .B(
        \pgld32[12] ), .C(\pgld16[12] ), .D(ph_word16_h) );
    snl_xnor2x0 \CONS/U195  ( .ZN(\CONS/n676 ), .A(\pk_pc_h[1] ), .B(
        \pk_pcs2_h[1] ) );
    snl_ao112x1 \PDOSEL/U46  ( .Z(PDLOUT[31]), .A(CDIN[31]), .B(\PDOSEL/n119 ), 
        .C(\ph_cpudout[31] ), .D(\pk_pdo_h[31] ) );
    snl_invx05 \CODEIF/U278  ( .ZN(\CODEIF/n3911 ), .A(\CODEIF/pfctr[15] ) );
    snl_nand02x1 \CODEIF/U344  ( .ZN(\CODEIF/n3880 ), .A(\CODEIF/pgctrinc[4] ), 
        .B(\CODEIF/n3945 ) );
    snl_invx05 \LDIS/U212  ( .ZN(\LDIS/n3136 ), .A(LIN[24]) );
    snl_nand02x1 \ALUIS/U174  ( .ZN(\ALUIS/n3668 ), .A(\pk_ada_h[10] ), .B(
        po_arsel_h) );
    snl_and02x1 \REG_2/U158  ( .Z(\ph_cpudout[28] ), .A(\ph_segset_h[28] ), 
        .B(seg_cnfg_h) );
    snl_nor02x1 \BLU/U333  ( .ZN(\BLU/n1472 ), .A(\BLU/n1548 ), .B(\BLU/n1547 
        ) );
    snl_xnor2x0 \CONS/U209  ( .ZN(\CONS/n693 ), .A(\pk_pc_h[14] ), .B(
        \pk_pcs1_h[14] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[15]  ( .Q(\ph_segset_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[15]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_oai222x0 \REGF/U584  ( .ZN(\REGF/RI_ACC[17] ), .A(\REGF/n8097 ), .B(
        \REGF/n8215 ), .C(\REGF/n8098 ), .D(\REGF/n8216 ), .E(\REGF/n8099 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U693  ( .ZN(\REGF/n8090 ), .A(PDLIN[20]) );
    snl_invx05 \REGF/U724  ( .ZN(\REGF/n8060 ), .A(\pgldi[30] ) );
    snl_oai122x0 \ADOSEL/U23  ( .ZN(\pgmuxout[12] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4125 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4126 ), .E(
        \ADOSEL/n4127 ) );
    snl_ffqrnx1 \MAIN/sprw_tap1_reg  ( .Q(\MAIN/sprw_tap1 ), .D(
        \pk_rwrit_h[65] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[11]  ( .Q(\pgld32[11] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexcl[11] ), .SE(lo_data_lth), .CP(SCLK
        ) );
    snl_nand02x1 \PDOSEL/U135  ( .ZN(\PDOSEL/n138 ), .A(\PDOSEL/n119 ), .B(
        CDIN[9]) );
    snl_and08x1 \CONS/U139  ( .Z(\CONS/n644 ), .A(\CONS/n692 ), .B(\CONS/n693 
        ), .C(\CONS/n694 ), .D(\CONS/n695 ), .E(\CONS/n696 ), .F(\CONS/n697 ), 
        .G(\CONS/n698 ), .H(\CONS/n691 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[26]  ( .Q(\ph_segset_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[26]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_nor02x1 \PDOSEL/U112  ( .ZN(\PDOSEL/n133 ), .A(\ph_cpudout[4] ), .B(
        \pk_pdo_h[4] ) );
    snl_invx05 \REGF/U703  ( .ZN(\REGF/n8105 ), .A(PDLIN[15]) );
    snl_oa112x1 \LBUS/U669  ( .Z(ph_d20lth), .A(\LBUS/n1450 ), .B(\LBUS/n1592 
        ), .C(\LBUS/n1417 ), .D(ph_timouth) );
    snl_nor02x2 \REGF/U392  ( .ZN(\REGF/n8228 ), .A(\ph_pdis_h[8] ), .B(
        \ph_pdis_h[7] ) );
    snl_ao022x1 \REGF/U433  ( .Z(\REGF/RI_PCOH[0] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[0]), .C(\stream4[32] ), .D(\REGF/n8053 ) );
    snl_aoi012x1 \ALUIS/U96  ( .ZN(\ALUIS/n3751 ), .A(\pgldi[30] ), .B(srcbsel
        ), .C(allfbsel) );
    snl_oai112x0 \LBUS/U559  ( .ZN(\LBUS/temp1[2] ), .A(\LBUS/n1395 ), .B(
        \LBUS/n1396 ), .C(\LBUS/n1397 ), .D(\LBUS/n1398 ) );
    snl_muxi21x1 \BLU/U439  ( .ZN(\BLU/n1579 ), .A(\BLU/n1576 ), .B(
        \BLU/n1575 ), .S(\poalufnc[1] ) );
    snl_oai222x0 \REGF/U434  ( .ZN(\REGF/RI_EACC[31] ), .A(\REGF/n8054 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8057 ), .E(\REGF/n8058 ), 
        .F(\REGF/n8059 ) );
    snl_ao022x1 \REGF/U498  ( .Z(\REGF/RI_PCOL[27] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[27]), .C(\stream4[27] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U508  ( .Z(\REGF/RI_PCOL[17] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[17]), .C(\stream4[17] ), .D(\REGF/n8209 ) );
    snl_oai022x1 \REGF/U638  ( .ZN(\REGF/RI_TBAI[20] ), .A(\REGF/n8225 ), .B(
        \REGF/n8157 ), .C(\REGF/n8226 ), .D(\REGF/n8158 ) );
    snl_nand02x1 \ADOSEL/U88  ( .ZN(\ADOSEL/n4154 ), .A(\pgbluext[31] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \CODEIF/U343  ( .ZN(\CODEIF/n3883 ), .A(\CODEIF/pgctrinc[5] ), 
        .B(\CODEIF/n3945 ) );
    snl_nand02x1 \ALUIS/U173  ( .ZN(\ALUIS/n3669 ), .A(\pk_ada_h[11] ), .B(
        po_arsel_h) );
    snl_nor04x0 \BLU/U334  ( .ZN(\BLU/n1475 ), .A(\BLU/n1546 ), .B(\BLU/n1548 
        ), .C(\BLU/n1549 ), .D(\BLU/n1545 ) );
    snl_ao022x1 \LDIS/U125  ( .Z(\pgld16[13] ), .A(ph_selldl), .B(\pgld32[13] 
        ), .C(ph_selldh), .D(\pgld32[29] ) );
    snl_invx05 \LDIS/U215  ( .ZN(\LDIS/n3161 ), .A(LIN[10]) );
    snl_xor2x0 \LDCHK/U59  ( .Z(\LDCHK/n3259 ), .A(\LDCHK/n3284 ), .B(
        \LDCHK/n3285 ) );
    snl_xnor2x0 \CONS/U192  ( .ZN(\CONS/n673 ), .A(\pgsdprlh[19] ), .B(
        \CONS/SACO[15] ) );
    snl_oai012x1 \PDOSEL/U41  ( .ZN(PDH[57]), .A(\PDOSEL/n111 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_ao022x1 \LDIS/U102  ( .Z(\pgldi[2] ), .A(ph_word32_h), .B(\pgld32[2] ), 
        .C(\pgld16[2] ), .D(ph_word16_h) );
    snl_nand12x1 \CMPX/U13  ( .ZN(ph_lbslock_h), .A(lbus_locken_h), .B(
        \CMPX/n1048 ) );
    snl_ao112x1 \PDOSEL/U66  ( .Z(PDLOUT[29]), .A(CDIN[29]), .B(\PDOSEL/n119 ), 
        .C(\ph_cpudout[29] ), .D(\pk_pdo_h[29] ) );
    snl_xor2x0 \CODEIF/U364  ( .Z(\CODEIF/n3939 ), .A(CDOUT[30]), .B(
        \CODEIF/n4024 ) );
    snl_nand02x1 \ALUIS/U154  ( .ZN(\ALUIS/n3687 ), .A(\pk_ada_h[29] ), .B(
        po_arsel_h) );
    snl_ao022x1 \BLUOS/U24  ( .Z(\pgbluext[5] ), .A(\pkbludgh[5] ), .B(
        ph_bit_h), .C(\pkdptout[5] ), .D(ph_word16_h) );
    snl_and08x1 \CONS/U30  ( .Z(ph_iyco_h), .A(\CONS/n520 ), .B(\CONS/n521 ), 
        .C(\CONS/n522 ), .D(\CONS/n523 ), .E(\CONS/n524 ), .F(\CONS/n525 ), 
        .G(\CONS/n526 ), .H(\CONS/n527 ) );
    snl_oai022x1 \BLU/U313  ( .ZN(\pkbludgh[3] ), .A(\BLU/n1464 ), .B(
        \BLU/n1501 ), .C(\BLU/n1502 ), .D(\BLU/n1503 ) );
    snl_oai222x0 \REGF/U583  ( .ZN(\REGF/RI_ACC[18] ), .A(\REGF/n8094 ), .B(
        \REGF/n8215 ), .C(\REGF/n8095 ), .D(\REGF/n8216 ), .E(\REGF/n8096 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U694  ( .ZN(\REGF/n8169 ), .A(\pgregadrh[19] ) );
    snl_invx05 \REGF/U704  ( .ZN(\REGF/n8179 ), .A(\pgregadrh[14] ) );
    snl_invx05 \CODEIF/U258  ( .ZN(\CODEIF/n3887 ), .A(\CODEIF/pfctr[7] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[17]  ( .Q(\ph_segset_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[17]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_aoi022x1 \ALUIS/U91  ( .ZN(\ALUIS/n3698 ), .A(\stream4[4] ), .B(
        immbsel), .C(\pk_adb_h[4] ), .D(po_brsel_h) );
    snl_xnor2x0 \CONS/U229  ( .ZN(\CONS/n528 ), .A(\pk_idcz_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[24]  ( .Q(\ph_segset_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[24]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_invx05 \REGF/U723  ( .ZN(\REGF/n8054 ), .A(\pgldi[31] ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[13]  ( .Q(\pgld32[13] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexcl[13] ), .SE(lo_data_lth), .CP(SCLK
        ) );
    snl_oai023x0 \CONS/U119  ( .ZN(\CONS/n637 ), .A(\CONS/n638 ), .B(
        ph_wrdsrc_h), .C(\pk_saseo_h[0] ), .D(\CONS/n542 ), .E(\CONS/n548 ) );
    snl_nor02x1 \PDOSEL/U115  ( .ZN(\PDOSEL/n135 ), .A(\ph_cpudout[27] ), .B(
        \pk_pdo_h[27] ) );
    snl_nor02x1 \LBUS/U649  ( .ZN(\LBUS/n1604 ), .A(\LBUS/n1601 ), .B(
        \LBUS/n1458 ) );
    snl_oai122x0 \ADOSEL/U24  ( .ZN(\pgmuxout[13] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4128 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4129 ), .E(
        \ADOSEL/n4130 ) );
    snl_muxi21x1 \LDIS/U189  ( .ZN(\LDIS/ldexch[21] ), .A(\LDIS/n3142 ), .B(
        \LDIS/n3141 ), .S(\LDIS/n3165 ) );
    snl_nor02x1 \PDOSEL/U132  ( .ZN(\PDOSEL/n127 ), .A(\ph_cpudout[11] ), .B(
        \pk_pdo_h[11] ) );
    snl_ao022x1 \REGF/U413  ( .Z(\REGF/RI_PCOH[20] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[20]), .C(\stream4[52] ), .D(\REGF/n8053 ) );
    snl_aoi013x0 \LBUS/U579  ( .ZN(ph_stdatlth), .A(\LBUS/n1430 ), .B(LDS), 
        .C(\LBUS/n1440 ), .D(\LBUS/n1441 ) );
    snl_nand02x2 \REGF/U377  ( .ZN(\REGF/n8055 ), .A(po_ldis_h), .B(
        \REGF/n8059 ) );
    snl_or08x1 \REGF/U656  ( .Z(pk_excp_h), .A(\REGF/RO_PSTA[19] ), .B(
        \REGF/RO_PSTA[20] ), .C(\REGF/RO_PSTA[17] ), .D(\REGF/RO_PSTA[18] ), 
        .E(\REGF/RO_PSTA[22] ), .F(CDOUT[59]), .G(\REGF/RO_PSTA[21] ), .H(
        \REGF/RO_PSTA[16] ) );
    snl_and02x1 \REGF/U828  ( .Z(\REGF/n8222 ), .A(\REGF/n8223 ), .B(
        \REGF/n8232 ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[8]  ( .Q(\REGF/RO_LLPSAS[10] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[8] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_and02x1 \ALUIS/U8  ( .Z(\ALUIS/n3641 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3668 ) );
    snl_ao022x1 \LDIS/U99  ( .Z(\pgld16[0] ), .A(ph_selldl), .B(\pgld32[0] ), 
        .C(ph_selldh), .D(\pgld32[16] ) );
    snl_nor02x1 \LBUS/U627  ( .ZN(\LBUS/n1598 ), .A(\LBUS/n1452 ), .B(
        \LBUS/ilt[0] ) );
    snl_invx05 \BLU/U398  ( .ZN(\BLU/n1482 ), .A(\pgld16[10] ) );
    snl_invx05 \BLU/U419  ( .ZN(\BLU/n1551 ), .A(\BLU/n1501 ) );
    snl_and08x1 \CONS/U150  ( .Z(\CONS/n527 ), .A(\CONS/n715 ), .B(\CONS/n716 
        ), .C(\CONS/n717 ), .D(\CONS/n718 ), .E(\CONS/n719 ), .F(\CONS/n720 ), 
        .G(\CONS/n721 ), .H(\CONS/n714 ) );
    snl_ao022x1 \REG_2/U131  ( .Z(\ph_cpudout[1] ), .A(\ph_segset_h[1] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[1] ), .D(ret_cont_h) );
    snl_invx05 \PDOSEL/U83  ( .ZN(\PDOSEL/n80 ), .A(CDIN[36]) );
    snl_ao222x1 \CODEIF/U211  ( .Z(\CODEIF/n3858 ), .A(PA[20]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[17] ), .E(cif_byte), .F(PDLIN[17]
        ) );
    snl_xnor2x0 \CODEIF/U381  ( .ZN(\CODEIF/n3976 ), .A(CPIN[2]), .B(CDIN[37])
         );
    snl_xor2x0 \CODEIF/U400  ( .Z(\CODEIF/n3961 ), .A(\CODEIF/n3957 ), .B(
        \CODEIF/n4036 ) );
    snl_xnor2x0 \CONS/U260  ( .ZN(\CONS/n348 ), .A(\pk_idcx_h[3] ), .B(
        \pk_indx_h[3] ) );
    snl_oai122x0 \CODEIF/U236  ( .ZN(\CODEIF/pfctr415[15] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3911 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3912 ), .E(
        \CODEIF/n3913 ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[3]  ( .Q(\pgld32[3] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[3] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_aoi012x1 \LBUS/U600  ( .ZN(\LBUS/n1421 ), .A(stage_b), .B(\LBUS/n1438 
        ), .C(word32odtrh) );
    snl_xnor2x0 \CONS/U247  ( .ZN(\CONS/n730 ), .A(\pk_idcx_h[22] ), .B(
        \pk_indx_h[22] ) );
    snl_xnor2x0 \CONS/U177  ( .ZN(\CONS/n654 ), .A(\pgsdprlh[10] ), .B(
        \pk_saco_lh[10] ) );
    snl_nand02x1 \ALUIS/U53  ( .ZN(\pgaluinb[5] ), .A(\ALUIS/n3700 ), .B(
        \ALUIS/n3701 ) );
    snl_oai222x2 \REGF/U389  ( .ZN(\REGF/RI_SRA12M[27] ), .A(\REGF/n8054 ), 
        .B(\REGF/n8051 ), .C(\REGF/n8227 ), .D(\REGF/n8153 ), .E(\REGF/n8228 ), 
        .F(\REGF/n8058 ) );
    snl_oai222x0 \REGF/U441  ( .ZN(\REGF/RI_EACC[24] ), .A(\REGF/n8076 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8077 ), .E(\REGF/n8078 ), 
        .F(\REGF/n8059 ) );
    snl_ao2222x1 \REGF/U541  ( .Z(\REGF/RI_SRDA[16] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[16]), .C(\pgldi[16] ), .D(\REGF/n8210 ), .E(\stream3[16] ), .F(
        \REGF/n8211 ), .G(\pkdptout[16] ), .H(\REGF/n8212 ) );
    snl_and02x1 \REGF/U566  ( .Z(\REGF/RO_LPSAS2156[8] ), .A(ph_sastlth), .B(
        \REGF/RO_PSTA[21] ) );
    snl_nand02x1 \ADOSEL/U112  ( .ZN(\ADOSEL/n4091 ), .A(\pgbluext[16] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U74  ( .ZN(\pgaluinb[26] ), .A(\ALUIS/n3742 ), .B(
        \ALUIS/n3743 ) );
    snl_invx05 \REGF/U671  ( .ZN(\REGF/n8126 ), .A(PDLIN[8]) );
    snl_nand02x1 \MAIN/U122  ( .ZN(\MAIN/*cell*4603/U10/CONTROL1 ), .A(
        \MAIN/n3613 ), .B(\MAIN/n3614 ) );
    snl_nor02x1 \LDCHK/U37  ( .ZN(\LDCHK/n3245 ), .A(\LDCHK/n3240 ), .B(
        \LDCHK/n3246 ) );
    snl_mux21x1 \ALUSHT/U38  ( .Z(\pkdptout[14] ), .A(\ALUSHT/pkshtout[14] ), 
        .B(\ALUSHT/pkaluout[14] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U79  ( .Z(\CONS/n597 ), .A(\pk_pcs1_h[3] ), .B(
        \pk_pc_h[3] ) );
    snl_invx05 \REGF/U771  ( .ZN(\REGF/n8174 ), .A(\pgsdprlh[17] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[1]  ( .Q(\REGF/RO_LLPSAS[1] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[1] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_nand02x1 \ADOSEL/U109  ( .ZN(\ADOSEL/n4127 ), .A(\pgbluext[28] ), .B(
        \ADOSEL/n4156 ) );
    snl_ao222x1 \CODEIF/U196  ( .Z(\CODEIF/n3843 ), .A(PA[5]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[2] ), .E(cif_byte), .F(PDLIN[2])
         );
    snl_and02x1 \MAIN/U139  ( .Z(ph_ltwt_h), .A(ph_filewr_h), .B(ltffsel) );
    snl_invx05 \LDIS/U150  ( .ZN(\LDIS/n3121 ), .A(\pgld32[21] ) );
    snl_mux21x1 \ALUSHT/U23  ( .Z(\pkdptout[28] ), .A(\ALUSHT/pkshtout[28] ), 
        .B(\ALUSHT/pkaluout[28] ), .S(\ALUSHT/n3112 ) );
    snl_invx05 \LBUS/U690  ( .ZN(\LBUS/n_2439 ), .A(\LBUS/n1399 ) );
    snl_xor2x0 \CONS/U62  ( .Z(\CONS/n579 ), .A(\CONS/SACO[10] ), .B(
        \pgsdprlh[14] ) );
    snl_oai022x1 \SAEXE/U107  ( .ZN(ph_lwdsrch), .A(\SAEXE/n413 ), .B(
        \SAEXE/n418 ), .C(\SAEXE/n415 ), .D(\SAEXE/n419 ) );
    snl_xor2x0 \CODEIF/U336  ( .Z(\CODEIF/n4019 ), .A(CDOUT[6]), .B(
        \CODEIF/n4018 ) );
    snl_aoi012x1 \ALUIS/U106  ( .ZN(\ALUIS/n3743 ), .A(\pgldi[26] ), .B(
        srcbsel), .C(allfbsel) );
    snl_invx05 \LDCHK/U123  ( .ZN(\LDCHK/n3312 ), .A(\LDCHK/n3296 ) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[6]  ( .Q(\REG_2/ph_retcnt_h[6] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[6]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_oai012x1 \PDOSEL/U34  ( .ZN(PDH[50]), .A(\PDOSEL/n104 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_invx05 \BLU/U341  ( .ZN(\BLU/n1523 ), .A(\poalufnc[0] ) );
    snl_invx05 \CODEIF/U281  ( .ZN(\CODEIF/n3909 ), .A(PDLIN[14]) );
    snl_xnor2x0 \LDCHK/U104  ( .ZN(\LDCHK/n3281 ), .A(\pgmuxout[27] ), .B(
        \pgmuxout[28] ) );
    snl_and34x0 \LBUS/U587  ( .Z(ph_bdstenh), .A(ph_btsrdaselh), .B(LRQ), .C(
        \LBUS/n1441 ), .D(ph_bit_h) );
    snl_nand03x0 \BLU/U366  ( .ZN(\BLU/n1550 ), .A(\BLU/n1483 ), .B(
        \BLU/n1486 ), .C(\BLU/n1480 ) );
    snl_xor2x0 \CODEIF/U311  ( .Z(\CODEIF/n3982 ), .A(\CODEIF/n3983 ), .B(
        \CODEIF/n3984 ) );
    snl_nand02x1 \ALUIS/U48  ( .ZN(\pgaluinb[0] ), .A(\ALUIS/n3690 ), .B(
        \ALUIS/n3691 ) );
    snl_aoi022x1 \ALUIS/U121  ( .ZN(\ALUIS/n3692 ), .A(\stream4[1] ), .B(
        immbsel), .C(\pk_adb_h[1] ), .D(po_brsel_h) );
    snl_invx05 \ADOSEL/U76  ( .ZN(\ADOSEL/n4119 ), .A(\pkdptout[26] ) );
    snl_muxi21x1 \LDIS/U177  ( .ZN(\LDIS/ldexcl[10] ), .A(\LDIS/n3161 ), .B(
        \LDIS/n3162 ), .S(\LDIS/n3134 ) );
    snl_or08x1 \CONS/U45  ( .Z(\CONS/n559 ), .A(\CONS/n560 ), .B(\CONS/n561 ), 
        .C(\CONS/n562 ), .D(\CONS/n563 ), .E(\CONS/n564 ), .F(\CONS/n565 ), 
        .G(\CONS/n566 ), .H(\CONS/n567 ) );
    snl_nand02x1 \SAEXE/U120  ( .ZN(\SAEXE/n427 ), .A(\SAEXE/n411 ), .B(
        \SAEXE/n429 ) );
    snl_ffqrnx1 \LBUS/ilt_reg[2]  ( .Q(\LBUS/ilt[2] ), .D(\LBUS/temp1[2] ), 
        .RN(n10734), .CP(SCLK) );
    snl_nand12x2 \PDOSEL/U13  ( .ZN(\PDOSEL/n75 ), .A(\PDOSEL/n223 ), .B(
        code_area_h) );
    snl_nand02x1 \PDOSEL/U160  ( .ZN(\PDOSEL/n136 ), .A(CDIN[12]), .B(
        \PDOSEL/n119 ) );
    snl_oai022x1 \REGF/U466  ( .ZN(\REGF/RI_DPR[27] ), .A(\REGF/n8058 ), .B(
        \REGF/n8151 ), .C(\REGF/n8152 ), .D(\REGF/n8153 ) );
    snl_muxi21x1 \REGF/U833  ( .ZN(\REGF/n8213 ), .A(\REGF/n8244 ), .B(PDLIN
        [0]), .S(\ph_pdis_h[9] ) );
    snl_oai222x0 \REGF/U598  ( .ZN(\REGF/RI_ACC[3] ), .A(\REGF/n8139 ), .B(
        \REGF/n8215 ), .C(\REGF/n8140 ), .D(\REGF/n8216 ), .E(\REGF/n8141 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U756  ( .ZN(\REGF/n8196 ), .A(\pgsdprlh[6] ) );
    snl_invx05 \REGF/U814  ( .ZN(\REGF/n8149 ), .A(\pkdptout[0] ) );
    snl_invx05 \ADOSEL/U51  ( .ZN(\ADOSEL/n4111 ), .A(\pkdptout[7] ) );
    snl_invx05 \PDOSEL/U98  ( .ZN(\PDOSEL/n102 ), .A(CDIN[48]) );
    snl_nand02x1 \PDOSEL/U147  ( .ZN(\PDOSEL/n164 ), .A(CDIN[23]), .B(
        \PDOSEL/n119 ) );
    snl_xor2x0 \LDCHK/U80  ( .Z(\LDCHK/n3269 ), .A(\LDCHK/n3305 ), .B(
        \LDCHK/n3306 ) );
    snl_invx05 \CODEIF/U264  ( .ZN(\CODEIF/n3878 ), .A(\CODEIF/pfctr[4] ) );
    snl_xnor2x0 \CONS/U215  ( .ZN(\CONS/n700 ), .A(\pk_pc_h[8] ), .B(
        \pk_pcs1_h[8] ) );
    snl_nand02x1 \BLU/U383  ( .ZN(\BLU/n1504 ), .A(\BLU/n1568 ), .B(
        \BLU/n1561 ) );
    snl_nor02x1 \BLU/U402  ( .ZN(\BLU/n1573 ), .A(accasel), .B(all0asel) );
    snl_nand23x1 \LBUS/U562  ( .ZN(ph_lberr), .A(\LBUS/n1402 ), .B(
        \LBUS/lnsa_err ), .C(\LBUS/n1403 ) );
    snl_and02x1 \REG_2/U144  ( .Z(\ph_cpudout[14] ), .A(\ph_segset_h[14] ), 
        .B(seg_cnfg_h) );
    snl_ao022x1 \REGF/U408  ( .Z(\REGF/RI_PCOH[25] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[25]), .C(\stream4[57] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U453  ( .ZN(\REGF/RI_EACC[12] ), .A(\REGF/n8112 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8113 ), .E(\REGF/n8114 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U483  ( .ZN(\REGF/RI_DPR[10] ), .A(\REGF/n8187 ), .B(
        \REGF/n8160 ), .C(\REGF/n8188 ), .D(\REGF/n8162 ), .E(\REGF/n8120 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U513  ( .Z(\REGF/RI_PCOL[12] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[12]), .C(\stream4[12] ), .D(\REGF/n8209 ) );
    snl_invx05 \REGF/U738  ( .ZN(\REGF/n8082 ), .A(\pgldi[22] ) );
    snl_muxi21x1 \LDIS/U192  ( .ZN(\LDIS/ldexch[18] ), .A(\LDIS/n3148 ), .B(
        \LDIS/n3147 ), .S(\LDIS/n3165 ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[24]  ( .Q(\pgld32[24] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[24] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[17]  ( .Q(\pgld32[17] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[17] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_nor03x0 \CONS/U125  ( .ZN(\CONS/n656 ), .A(\CONS/n573 ), .B(
        \CONS/n571 ), .C(\CONS/n572 ) );
    snl_nor02x1 \PDOSEL/U129  ( .ZN(\PDOSEL/n143 ), .A(\pk_pdo_h[14] ), .B(
        \ph_cpudout[14] ) );
    snl_oai122x0 \ADOSEL/U18  ( .ZN(\pgmuxout[7] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4110 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4111 ), .E(
        \ADOSEL/n4112 ) );
    snl_oa023x1 \LBUS/U652  ( .Z(\LBUS/n1603 ), .A(LRQ), .B(\LBUS/ilt[4] ), 
        .C(\LBUS/n1455 ), .D(\LBUS/n1461 ), .E(ph_timouth) );
    snl_xor2x0 \CODEIF/U243  ( .Z(\CODEIF/n3930 ), .A(\CODEIF/n3931 ), .B(
        \CODEIF/n3932 ) );
    snl_invx05 \LBUS/U675  ( .ZN(\LBUS/n1423 ), .A(\LBUS/n1600 ) );
    snl_xor2x0 \CONS/U87  ( .Z(\CONS/n605 ), .A(\pk_idcz_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_xor2x0 \CONS/U102  ( .Z(\CONS/n620 ), .A(\pk_idcx_h[4] ), .B(
        \pk_indx_h[4] ) );
    snl_xnor2x0 \CONS/U232  ( .ZN(\CONS/n718 ), .A(\pk_idcy_h[16] ), .B(
        \pk_indy_h[16] ) );
    snl_invx05 \BLU/U425  ( .ZN(\BLU/n1531 ), .A(\BLU/n1477 ) );
    snl_oai222x0 \REGF/U491  ( .ZN(\REGF/RI_DPR[2] ), .A(\REGF/n8203 ), .B(
        \REGF/n8160 ), .C(\REGF/n8204 ), .D(\REGF/n8162 ), .E(\REGF/n8144 ), 
        .F(\REGF/n8151 ) );
    snl_ao2222x1 \REGF/U534  ( .Z(\REGF/RI_SRDA[23] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[23]), .C(\pgldi[23] ), .D(\REGF/n8210 ), .E(\stream3[23] ), .F(
        \REGF/n8211 ), .G(\pkdptout[23] ), .H(\REGF/n8212 ) );
    snl_oai022x1 \REGF/U604  ( .ZN(\REGF/RI_SPR[25] ), .A(\REGF/n8155 ), .B(
        \REGF/n8218 ), .C(\REGF/n8219 ), .D(\REGF/n8156 ) );
    snl_oai222x0 \REGF/U623  ( .ZN(\REGF/RI_SPR[6] ), .A(\REGF/n8195 ), .B(
        \REGF/n8220 ), .C(\REGF/n8196 ), .D(\REGF/n8221 ), .E(\REGF/n8132 ), 
        .F(\REGF/n8218 ) );
    snl_invx1 \ALUIS/U26  ( .ZN(\pgaluina[1] ), .A(\ALUIS/n3653 ) );
    snl_and02x1 \LDIS/U229  ( .Z(\LDIS/n3165 ), .A(\pgsadrh[0] ), .B(
        ph_word32_h) );
    snl_xor2x0 \LDCHK/U65  ( .Z(\LDCHK/n3295 ), .A(\pgld32[4] ), .B(
        \LDCHK/n3294 ) );
    snl_oai022x1 \BLU/U308  ( .ZN(\pkbludgh[8] ), .A(\BLU/n1464 ), .B(
        \BLU/n1486 ), .C(\BLU/n1487 ), .D(\BLU/n1488 ) );
    snl_invx05 \REGF/U794  ( .ZN(\REGF/n8066 ), .A(\pkdptout[28] ) );
    snl_ao022x1 \BLUOS/U18  ( .Z(\pgbluext[30] ), .A(\pkbludgh[14] ), .B(
        ph_bit_h), .C(\pkdptout[14] ), .D(ph_word16_h) );
    snl_invx05 \MAIN/U170  ( .ZN(ph_stregwt_h), .A(\MAIN/n3616 ) );
    snl_ao022x1 \LDIS/U119  ( .Z(\pgld16[10] ), .A(ph_selldl), .B(\pgld32[10] 
        ), .C(ph_selldh), .D(\pgld32[26] ) );
    snl_nand02x1 \ADOSEL/U93  ( .ZN(\ADOSEL/n4150 ), .A(\pgbluext[27] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \MAIN/U157  ( .ZN(\MAIN/n3617 ), .A(pkaccovf), .B(st_exectl)
         );
    snl_invx05 \LDCHK/U42  ( .ZN(\LDCHK/n3255 ), .A(\pgld32[31] ) );
    snl_xnor2x0 \CONS/U189  ( .ZN(\CONS/n668 ), .A(\pgsdprlh[18] ), .B(
        \CONS/SACO[14] ) );
    snl_xor2x0 \CODEIF/U358  ( .Z(\CODEIF/n3932 ), .A(CDIN[58]), .B(
        \CODEIF/n3946 ) );
    snl_nand02x1 \ALUIS/U168  ( .ZN(\ALUIS/n3674 ), .A(\pk_ada_h[16] ), .B(
        po_arsel_h) );
    snl_ao022x1 \REGF/U501  ( .Z(\REGF/RI_PCOL[24] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[24]), .C(\stream4[24] ), .D(\REGF/n8209 ) );
    snl_ao2222x1 \REGF/U526  ( .Z(\REGF/RI_SRDA[31] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[31]), .C(\pgldi[31] ), .D(\REGF/n8210 ), .E(\stream3[31] ), .F(
        \REGF/n8211 ), .G(\pkdptout[31] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U616  ( .ZN(\REGF/RI_SPR[13] ), .A(\REGF/n8181 ), .B(
        \REGF/n8220 ), .C(\REGF/n8182 ), .D(\REGF/n8221 ), .E(\REGF/n8111 ), 
        .F(\REGF/n8218 ) );
    snl_and12x1 \REGF/U631  ( .Z(\REGF/RI_STAT[4] ), .A(\REGF/n8222 ), .B(
        PDLIN[30]) );
    snl_nand02x1 \ALUIS/U34  ( .ZN(\pgaluina[18] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3676 ) );
    snl_oai013x0 \MAIN/U162  ( .ZN(\MAIN/n3615 ), .A(baccsel), .B(po_cmfsel_h), 
        .C(po_opcsel_h), .D(ph_filewr_h) );
    snl_xor2x0 \LDCHK/U77  ( .Z(\LDCHK/n3265 ), .A(\LDCHK/n3303 ), .B(
        \LDCHK/n3304 ) );
    snl_aoi022x1 \CONS/U39  ( .ZN(\CONS/n544 ), .A(\CONS/n551 ), .B(
        \CONS/n546 ), .C(\pgsdprlh[4] ), .D(\pk_saco_lh[4] ) );
    snl_xor2x0 \LDCHK/U50  ( .Z(\LDCHK/n3268 ), .A(\LDCHK/n3269 ), .B(
        \LDCHK/n3270 ) );
    snl_invx05 \REGF/U786  ( .ZN(\REGF/n8131 ), .A(\pkdptout[6] ) );
    snl_nand02x1 \ADOSEL/U81  ( .ZN(\ADOSEL/n4118 ), .A(\pgbluext[9] ), .B(
        \ADOSEL/n4156 ) );
    snl_nor02x1 \MAIN/U145  ( .ZN(\MAIN/single_read ), .A(pgadrovfh), .B(
        \MAIN/n3631 ) );
    snl_oai112x0 \PDOSEL/U48  ( .ZN(PDLOUT[13]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n99 ), .C(\PDOSEL/n122 ), .D(\PDOSEL/n123 ) );
    snl_invx05 \REGF/U763  ( .ZN(\REGF/n8161 ), .A(\pgsdprlh[23] ) );
    snl_invx05 \ADOSEL/U64  ( .ZN(\ADOSEL/n4134 ), .A(\pkdptout[31] ) );
    snl_invx05 \CODEIF/U251  ( .ZN(\CODEIF/n3863 ), .A(write_pr_h) );
    snl_invx05 \CODEIF/U276  ( .ZN(\CODEIF/n3914 ), .A(\CODEIF/pfctr[16] ) );
    snl_invx1 \ALUIS/U13  ( .ZN(\pgaluina[0] ), .A(\ALUIS/n3645 ) );
    snl_and02x1 \REG_2/U156  ( .Z(\ph_cpudout[26] ), .A(\ph_segset_h[26] ), 
        .B(seg_cnfg_h) );
    snl_nand02x1 \BLU/U391  ( .ZN(\BLU/n1468 ), .A(\BLU/n1567 ), .B(
        \BLU/n1561 ) );
    snl_aoi012x1 \ALUIS/U98  ( .ZN(\ALUIS/n3695 ), .A(\pgldi[2] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_muxi21x1 \LDIS/U180  ( .ZN(\LDIS/ldexch[30] ), .A(\LDIS/n3154 ), .B(
        \LDIS/n3153 ), .S(\LDIS/n3165 ) );
    snl_nand12x1 \LBUS/U570  ( .ZN(\LBUS/*cell*3982/U201/CONTROL1 ), .A(
        \LBUS/*cell*3982/U119/CONTROL1 ), .B(\LBUS/n1400 ) );
    snl_xnor2x0 \CONS/U207  ( .ZN(\CONS/n698 ), .A(\pk_pc_h[11] ), .B(
        \pk_pcs1_h[11] ) );
    snl_nor02x1 \BLU/U410  ( .ZN(\BLU/n1583 ), .A(\BLU/n1556 ), .B(\BLU/n1558 
        ) );
    snl_nor04x0 \CONS/U137  ( .ZN(\CONS/n645 ), .A(\CONS/n686 ), .B(
        \CONS/n682 ), .C(\CONS/n589 ), .D(\CONS/n590 ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[7]  ( .Q(\pgld32[7] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[7] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_nor02x1 \LBUS/U640  ( .ZN(\LBUS/n1424 ), .A(word32odtrh), .B(
        ph_lbslock_h) );
    snl_invx05 \LBUS/U667  ( .ZN(\LBUS/n1407 ), .A(\LBUS/n1445 ) );
    snl_xor2x0 \CONS/U110  ( .Z(\CONS/n628 ), .A(\pk_idcw_h[8] ), .B(
        \pk_indw_h[8] ) );
    snl_xor2x0 \CONS/U95  ( .Z(\CONS/n613 ), .A(\pk_idcy_h[23] ), .B(
        \pk_indy_h[23] ) );
    snl_oai123x2 \LBUS/U557  ( .ZN(ph_lbend), .A(\LBUS/n1406 ), .B(
        \LBUS/n1407 ), .C(\LBUS/n1408 ), .D(\LBUS/n1407 ), .E(\LBUS/n1409 ), 
        .F(\LBUS/n1410 ) );
    snl_xnor2x0 \CONS/U220  ( .ZN(\CONS/n703 ), .A(\pk_idcz_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_muxi21x1 \BLU/U437  ( .ZN(\BLU/n1520 ), .A(\BLU/n1573 ), .B(
        \pk_stat_h[1] ), .S(eaccasel) );
    snl_or04x1 \REGF/U821  ( .Z(\REGF/n8243 ), .A(\REGF/RO_ACC[26] ), .B(
        \REGF/RO_ACC[25] ), .C(\REGF/RO_ACC[30] ), .D(pk_sign_h) );
    snl_mux21x1 \SHTCD/U12  ( .Z(\phshtd[5] ), .A(\pgld16[5] ), .B(
        \stream4[5] ), .S(immbsel) );
    snl_invx05 \LBUS/U609  ( .ZN(\LBUS/n1453 ), .A(\LBUS/ilt[5] ) );
    snl_oai222x0 \REGF/U474  ( .ZN(\REGF/RI_DPR[19] ), .A(\REGF/n8169 ), .B(
        \REGF/n8160 ), .C(\REGF/n8170 ), .D(\REGF/n8162 ), .E(\REGF/n8093 ), 
        .F(\REGF/n8151 ) );
    snl_invx05 \REGF/U806  ( .ZN(\REGF/n8098 ), .A(\pkdptout[17] ) );
    snl_aoi013x2 \CODEIF/U218  ( .ZN(pgperrh), .A(\CODEIF/n3923 ), .B(
        \CODEIF/n3924 ), .C(\CODEIF/n3925 ), .D(CROE) );
    snl_xnor2x0 \CODEIF/U388  ( .ZN(\CODEIF/n3984 ), .A(CDIN[21]), .B(CDIN[19]
        ) );
    snl_xnor2x0 \CODEIF/U409  ( .ZN(\CODEIF/n4039 ), .A(CDOUT[35]), .B(CDOUT
        [38]) );
    snl_and02x1 \REG_2/U138  ( .Z(\ph_cpudout[8] ), .A(\ph_segset_h[8] ), .B(
        seg_cnfg_h) );
    snl_xnor2x0 \CONS/U269  ( .ZN(\CONS/n749 ), .A(\pk_idcw_h[12] ), .B(
        \pk_indw_h[12] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[13]  ( .Q(\ph_segset_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[13]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_invx05 \REGF/U744  ( .ZN(\REGF/n8097 ), .A(\pgldi[17] ) );
    snl_nand02x1 \ADOSEL/U43  ( .ZN(\ADOSEL/n4155 ), .A(ph_word32_h), .B(
        \pgsadrh[0] ) );
    snl_ffqrnx1 \MAIN/astregw_tap1_reg  ( .Q(\MAIN/astregw_tap1 ), .D(
        \MAIN/*cell*4603/U14/CONTROL1 ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nand02x1 \PDOSEL/U155  ( .ZN(\PDOSEL/n152 ), .A(CDIN[17]), .B(
        \PDOSEL/n119 ) );
    snl_nor03x0 \CONS/U159  ( .ZN(\CONS/n341 ), .A(\CONS/n633 ), .B(
        \CONS/n631 ), .C(\CONS/n632 ) );
    snl_invx05 \LDCHK/U92  ( .ZN(\LDCHK/n3239 ), .A(\pgld32[27] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[20]  ( .Q(\ph_segset_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[20]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_oai2222x0 \REGF/U359  ( .ZN(\REGF/RI_SRA12M[15] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8105 ), .C(\REGF/n8103 ), .D(\REGF/n8051 ), .E(\REGF/n8177 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8178 ) );
    snl_invx05 \REGF/U678  ( .ZN(\REGF/n8154 ), .A(\pgsdprhh[30] ) );
    snl_mux21x1 \ALUSHT/U31  ( .Z(\pkdptout[20] ), .A(\ALUSHT/pkshtout[20] ), 
        .B(\ALUSHT/pkaluout[20] ), .S(\ALUSHT/n3112 ) );
    snl_invx05 \LBUS/U682  ( .ZN(\LBUS/n1397 ), .A(\LBUS/nlt[3] ) );
    snl_xor2x0 \CONS/U70  ( .Z(\CONS/n588 ), .A(\pk_pc_h[10] ), .B(
        \pk_pcs2_h[10] ) );
    snl_oai022x1 \SAEXE/U115  ( .ZN(ph_word16h), .A(\SAEXE/n413 ), .B(
        \SAEXE/n414 ), .C(\SAEXE/n415 ), .D(\SAEXE/n426 ) );
    snl_oai012x1 \LDIS/U142  ( .ZN(\pgldi[28] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3128 ), .C(\LDIS/n3115 ) );
    snl_oai012x1 \PDOSEL/U26  ( .ZN(PDH[42]), .A(\PDOSEL/n96 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_oai2222x0 \REGF/U365  ( .ZN(\REGF/RI_SRA12M[5] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8135 ), .C(\REGF/n8133 ), .D(\REGF/n8051 ), .E(\REGF/n8197 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8198 ) );
    snl_ao2222x1 \REGF/U548  ( .Z(\REGF/RI_SRDA[9] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[9]), .C(\REGF/n8210 ), .D(\pgldi[9] ), .E(\REGF/n8211 ), .F(
        \stream3[9] ), .G(\REGF/n8212 ), .H(\pkdptout[9] ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[30]  ( .Q(\pgld32[30] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[30] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[29]  ( .Q(\pgld32[29] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[29] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_oai222x0 \REGF/U574  ( .ZN(\REGF/RI_ACC[27] ), .A(\REGF/n8067 ), .B(
        \REGF/n8215 ), .C(\REGF/n8068 ), .D(\REGF/n8216 ), .E(\REGF/n8069 ), 
        .F(\REGF/n8217 ) );
    snl_oai022x1 \REGF/U644  ( .ZN(\REGF/RI_TBAI[13] ), .A(\REGF/n8225 ), .B(
        \REGF/n8099 ), .C(\REGF/n8226 ), .D(\REGF/n8173 ) );
    snl_ffqsnx1 \CODEIF/pgfpwel_reg  ( .Q(CRWE), .D(pgrstith), .SN(
        \CODEIF/n3861 ), .CP(SCLK) );
    snl_nor02x1 \BLU/U353  ( .ZN(\BLU/n1568 ), .A(\pgbitnoh[2] ), .B(
        \pgbitnoh[3] ) );
    snl_xor2x0 \CODEIF/U293  ( .Z(\CODEIF/n3952 ), .A(\CODEIF/n3953 ), .B(
        \CODEIF/n3954 ) );
    snl_xor2x0 \CODEIF/U303  ( .Z(\CODEIF/n3970 ), .A(CDIN[53]), .B(
        \CODEIF/n3969 ) );
    snl_xor2x0 \CODEIF/U324  ( .Z(\CODEIF/n4001 ), .A(\CODEIF/n4002 ), .B(
        \CODEIF/n4003 ) );
    snl_aoi012x1 \ALUIS/U114  ( .ZN(\ALUIS/n3735 ), .A(\pgldi[22] ), .B(
        srcbsel), .C(allfbsel) );
    snl_aoi022x1 \ALUIS/U133  ( .ZN(\ALUIS/n3718 ), .A(\stream4[14] ), .B(
        immbsel), .C(\pk_adb_h[14] ), .D(po_brsel_h) );
    snl_xnor2x0 \LDCHK/U116  ( .ZN(\LDCHK/n3293 ), .A(\pgmuxout[0] ), .B(
        \pgmuxout[1] ) );
    snl_and02x1 \LBUS/U595  ( .Z(ph_lbe1_h), .A(phsaerrh), .B(\LBUS/MMBSEL )
         );
    snl_invx05 \BLU/U374  ( .ZN(\BLU/n1497 ), .A(\pgld16[5] ) );
    snl_muxi21x1 \LDIS/U165  ( .ZN(\LDIS/ldexcl[7] ), .A(\LDIS/n3137 ), .B(
        \LDIS/n3138 ), .S(\LDIS/n3134 ) );
    snl_mux21x1 \ALUSHT/U16  ( .Z(\pkdptout[5] ), .A(\ALUSHT/pkshtout[5] ), 
        .B(\ALUSHT/pkaluout[5] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U57  ( .Z(\CONS/n561 ), .A(\pgsdprlh[20] ), .B(
        \CONS/SACO[16] ) );
    snl_nand13x1 \SAEXE/U132  ( .ZN(\SAEXE/n418 ), .A(\pk_psae_h[0] ), .B(
        \SAEXE/n429 ), .C(\pk_psae_h[1] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[30]  ( .Q(\ph_segset_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[30]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[29]  ( .Q(\ph_segset_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[29]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_nand02x1 \SAEXE/U129  ( .ZN(\SAEXE/n415 ), .A(\pk_psae_h[7] ), .B(
        ph_saexe_sth) );
    snl_invx05 \CODEIF/U288  ( .ZN(\CODEIF/n3896 ), .A(\CODEIF/pfctr[10] ) );
    snl_nor02x1 \CODEIF/U318  ( .ZN(\CODEIF/n3925 ), .A(\CODEIF/n3930 ), .B(
        \CODEIF/n3933 ) );
    snl_aoi012x1 \ALUIS/U128  ( .ZN(\ALUIS/n3723 ), .A(\pgldi[16] ), .B(
        srcbsel), .C(allfbsel) );
    snl_nand02x1 \ALUIS/U41  ( .ZN(\pgaluina[25] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3683 ) );
    snl_and02x1 \UPIF/U13  ( .Z(\ph_pdis_h[7] ), .A(\pk_rread_h[44] ), .B(
        \UPIF/n1046 ) );
    snl_oai2222x0 \REGF/U380  ( .ZN(\REGF/RI_SRA12M[14] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8108 ), .C(\REGF/n8106 ), .D(\REGF/n8051 ), .E(\REGF/n8179 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8180 ) );
    snl_ao022x1 \REGF/U426  ( .Z(\REGF/RI_PCOH[7] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[7]), .C(\stream4[39] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U448  ( .ZN(\REGF/RI_EACC[17] ), .A(\REGF/n8097 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8098 ), .E(\REGF/n8099 ), 
        .F(\REGF/n8059 ) );
    snl_ao2222x1 \REGF/U553  ( .Z(\REGF/RI_SRDA[4] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[4]), .C(\pgldi[4] ), .D(\REGF/n8210 ), .E(\stream3[4] ), .F(
        \REGF/n8211 ), .G(\pkdptout[4] ), .H(\REGF/n8212 ) );
    snl_nand02x1 \ADOSEL/U100  ( .ZN(\ADOSEL/n4143 ), .A(\pgbluext[4] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U66  ( .ZN(\pgaluinb[18] ), .A(\ALUIS/n3726 ), .B(
        \ALUIS/n3727 ) );
    snl_nor02x1 \BLU/U348  ( .ZN(\BLU/n1563 ), .A(\pgbitnoh[0] ), .B(
        \pgbitnoh[1] ) );
    snl_invx05 \REGF/U663  ( .ZN(\REGF/n8114 ), .A(PDLIN[12]) );
    snl_ao022x1 \MAIN/U130  ( .Z(ph_shelter_h), .A(po_shelter_h2), .B(
        \MAIN/n3624 ), .C(po_shelter_h1), .D(\MAIN/n3625 ) );
    snl_invx05 \LDIS/U159  ( .ZN(\LDIS/n3127 ), .A(\pgld32[27] ) );
    snl_invx05 \ADOSEL/U58  ( .ZN(\ADOSEL/n4098 ), .A(\pkdptout[19] ) );
    snl_invx05 \LDCHK/U89  ( .ZN(\LDCHK/n3273 ), .A(LPIN[1]) );
    snl_invx05 \LBUS/U635  ( .ZN(\LBUS/n1404 ), .A(word32odtrh) );
    snl_nor04x0 \CONS/U142  ( .ZN(\CONS/n642 ), .A(\CONS/n597 ), .B(
        \CONS/n598 ), .C(\CONS/n599 ), .D(\CONS/n600 ) );
    snl_invx05 \PDOSEL/U91  ( .ZN(\PDOSEL/n108 ), .A(CDIN[54]) );
    snl_ao222x1 \CODEIF/U203  ( .Z(\CODEIF/n3850 ), .A(PA[12]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[9] ), .E(cif_byte), .F(PDLIN[9])
         );
    snl_xnor2x0 \CODEIF/U393  ( .ZN(\CODEIF/n3987 ), .A(CDIN[10]), .B(CDIN[11]
        ) );
    snl_xor2x0 \CODEIF/U412  ( .Z(\CODEIF/n3938 ), .A(\CODEIF/n4007 ), .B(
        \CODEIF/n4040 ) );
    snl_xnor2x0 \CONS/U272  ( .ZN(\CONS/n343 ), .A(\pk_idcw_h[14] ), .B(
        \pk_indw_h[14] ) );
    snl_invx05 \REGF/U778  ( .ZN(\REGF/n8188 ), .A(\pgsdprlh[10] ) );
    snl_oai122x0 \CODEIF/U224  ( .ZN(\CODEIF/pfctr415[3] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3875 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3876 ), .E(
        \CODEIF/n3877 ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[20]  ( .Q(\pgld32[20] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[20] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_xnor2x0 \CONS/U255  ( .ZN(\CONS/n350 ), .A(\pk_idcx_h[9] ), .B(
        \pk_indx_h[9] ) );
    snl_nand12x1 \BLU/U442  ( .ZN(\BLU/n1581 ), .A(ebaccsel), .B(
        \pk_stat_h[0] ) );
    snl_nand04x0 \LBUS/U612  ( .ZN(\LBUS/n1462 ), .A(LASIN), .B(LGR), .C(
        \LBUS/access_en_h ), .D(\LBUS/n1425 ) );
    snl_nor02x1 \CONS/U165  ( .ZN(\CONS/n542 ), .A(\CONS/n549 ), .B(
        \CONS/n544 ) );
    snl_invx05 \REGF/U686  ( .ZN(\REGF/n8159 ), .A(\pgregadrh[23] ) );
    snl_aoi022x1 \ALUIS/U83  ( .ZN(\ALUIS/n3706 ), .A(\stream4[8] ), .B(
        immbsel), .C(\pk_adb_h[8] ), .D(po_brsel_h) );
    snl_invx05 \REGF/U716  ( .ZN(\REGF/n8124 ), .A(\pgldi[8] ) );
    snl_invx05 \REGF/U731  ( .ZN(\REGF/n8070 ), .A(\pgldi[26] ) );
    snl_oai122x0 \ADOSEL/U11  ( .ZN(\pgmuxout[0] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4088 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4090 ), .E(
        \ADOSEL/n4091 ) );
    snl_nor02x1 \PDOSEL/U107  ( .ZN(\PDOSEL/n139 ), .A(\ph_cpudout[9] ), .B(
        \pk_pdo_h[9] ) );
    snl_oai122x0 \ADOSEL/U36  ( .ZN(\pgmuxout[25] ), .A(\ADOSEL/n4117 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4116 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4148 ) );
    snl_nor02x1 \PDOSEL/U120  ( .ZN(\PDOSEL/n155 ), .A(\pk_pdo_h[22] ), .B(
        \ph_cpudout[22] ) );
    snl_nand02x2 \REGF/U401  ( .ZN(\REGF/n8160 ), .A(ph_sais_h), .B(
        \REGF/n8151 ) );
    snl_oai222x0 \REGF/U443  ( .ZN(\REGF/RI_EACC[22] ), .A(\REGF/n8082 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8083 ), .E(\REGF/n8084 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U464  ( .ZN(\REGF/RI_EACC[1] ), .A(\REGF/n8145 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8146 ), .E(\REGF/n8147 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U481  ( .ZN(\REGF/RI_DPR[12] ), .A(\REGF/n8183 ), .B(
        \REGF/n8160 ), .C(\REGF/n8184 ), .D(\REGF/n8162 ), .E(\REGF/n8114 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U511  ( .Z(\REGF/RI_PCOL[14] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[14]), .C(\stream4[14] ), .D(\REGF/n8209 ) );
    snl_ao2222x1 \REGF/U536  ( .Z(\REGF/RI_SRDA[21] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[21]), .C(\pgldi[21] ), .D(\REGF/n8210 ), .E(\stream3[21] ), .F(
        \REGF/n8211 ), .G(\pkdptout[21] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U591  ( .ZN(\REGF/RI_ACC[10] ), .A(\REGF/n8118 ), .B(
        \REGF/n8215 ), .C(\REGF/n8119 ), .D(\REGF/n8216 ), .E(\REGF/n8120 ), 
        .F(\REGF/n8217 ) );
    snl_oai222x0 \REGF/U606  ( .ZN(\REGF/RI_SPR[23] ), .A(\REGF/n8159 ), .B(
        \REGF/n8220 ), .C(\REGF/n8161 ), .D(\REGF/n8221 ), .E(\REGF/n8081 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U796  ( .ZN(\REGF/n8071 ), .A(\pkdptout[26] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[5]  ( .Q(\REGF/RO_LLPSAS[7] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[5] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_invx05 \LDIS/U207  ( .ZN(\LDIS/n3139 ), .A(LIN[6]) );
    snl_nand02x1 \ADOSEL/U91  ( .ZN(\ADOSEL/n4152 ), .A(\pgbluext[29] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \CODEIF/U351  ( .ZN(\CODEIF/n3913 ), .A(\CODEIF/pgctrinc[15] 
        ), .B(\CODEIF/n3945 ) );
    snl_nand02x1 \ALUIS/U161  ( .ZN(\ALUIS/n3680 ), .A(\pk_ada_h[22] ), .B(
        po_arsel_h) );
    snl_xor2x0 \CODEIF/U376  ( .Z(\CODEIF/n4031 ), .A(\CODEIF/n3966 ), .B(
        \CODEIF/n3970 ) );
    snl_nand02x1 \ALUIS/U146  ( .ZN(\ALUIS/n3665 ), .A(\pk_ada_h[7] ), .B(
        po_arsel_h) );
    snl_ao022x1 \LDIS/U110  ( .Z(\pgldi[6] ), .A(ph_word32_h), .B(\pgld32[6] ), 
        .C(\pgld16[6] ), .D(ph_word16_h) );
    snl_oai012x1 \LDIS/U137  ( .ZN(\pgldi[23] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3123 ), .C(\LDIS/n3115 ) );
    snl_ao022x1 \CMPX/U26  ( .Z(ph_dprtrs_h), .A(ph_dprsel2_h), .B(
        ph_saexe_sth), .C(po_dprtrs_h), .D(\CMPX/n1047 ) );
    snl_xnor2x0 \CONS/U180  ( .ZN(\CONS/n658 ), .A(\pgsdprlh[13] ), .B(
        \pk_saco_lh[13] ) );
    snl_nor02x1 \BLU/U326  ( .ZN(\BLU/n1496 ), .A(\BLU/n1537 ), .B(\BLU/n1536 
        ) );
    snl_oai112x0 \PDOSEL/U53  ( .ZN(PDLOUT[19]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n105 ), .C(\PDOSEL/n130 ), .D(\PDOSEL/n131 ) );
    snl_sffqenrnx1 \REG_2/ph_retcnt_h_reg[2]  ( .Q(\REG_2/ph_retcnt_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[2]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_oai112x0 \PDOSEL/U74  ( .ZN(PDLOUT[8]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n94 ), .C(\PDOSEL/n180 ), .D(\PDOSEL/n181 ) );
    snl_invx05 \LDIS/U220  ( .ZN(\LDIS/n3158 ), .A(LIN[28]) );
    snl_oai022x1 \BLU/U301  ( .ZN(\pkbludgh[15] ), .A(\BLU/n1464 ), .B(
        \BLU/n1465 ), .C(\BLU/n1466 ), .D(\BLU/n1467 ) );
    snl_oai012x1 \MAIN/U155  ( .ZN(\MAIN/n3612 ), .A(\MAIN/ovferlth ), .B(
        st_exectl), .C(\MAIN/n3623 ) );
    snl_oai112x0 \PDOSEL/U58  ( .ZN(PDLOUT[26]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n112 ), .C(\PDOSEL/n140 ), .D(\PDOSEL/n141 ) );
    snl_xnor2x0 \LDCHK/U40  ( .ZN(\LDCHK/n3253 ), .A(\pgld32[16] ), .B(
        \LDCHK/n3254 ) );
    snl_nand02x2 \ALUIS/U24  ( .ZN(\pgaluina[4] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3662 ) );
    snl_oai222x0 \REGF/U621  ( .ZN(\REGF/RI_SPR[8] ), .A(\REGF/n8191 ), .B(
        \REGF/n8220 ), .C(\REGF/n8192 ), .D(\REGF/n8221 ), .E(\REGF/n8126 ), 
        .F(\REGF/n8218 ) );
    snl_oai022x1 \MAIN/U172  ( .ZN(\MAIN/n3625 ), .A(\MAIN/b_exec_stage ), .B(
        ph_dec_ch), .C(\MAIN/d_exec_stage ), .D(ph_dec_ah) );
    snl_xor2x0 \LDCHK/U67  ( .Z(\LDCHK/n3297 ), .A(\pgld32[1] ), .B(
        \pgld32[6] ) );
    snl_nor04x0 \REGF/U816  ( .ZN(\REGF/n8239 ), .A(\REGF/n8240 ), .B(
        \REGF/n8241 ), .C(\REGF/n8242 ), .D(\REGF/n8243 ) );
    snl_nor02x1 \CODEIF/U241  ( .ZN(\CODEIF/n3926 ), .A(\CODEIF/wprotect0 ), 
        .B(\CODEIF/n3927 ) );
    snl_invx05 \LBUS/U677  ( .ZN(\LBUS/n1409 ), .A(\LBUS/n1598 ) );
    snl_and08x1 \CONS/U29  ( .Z(ph_ixco_h), .A(\CONS/n346 ), .B(\CONS/n347 ), 
        .C(\CONS/n348 ), .D(\CONS/n349 ), .E(\CONS/n350 ), .F(\CONS/n351 ), 
        .G(\CONS/n518 ), .H(\CONS/n519 ) );
    snl_xor2x0 \CONS/U85  ( .Z(\CONS/n603 ), .A(\pk_idcz_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_xor2x0 \CONS/U100  ( .Z(\CONS/n618 ), .A(\pk_idcy_h[15] ), .B(
        \pk_indy_h[15] ) );
    snl_xnor2x0 \CONS/U230  ( .ZN(\CONS/n530 ), .A(\pk_idcz_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_and02x1 \REG_2/U161  ( .Z(\ph_cpudout[31] ), .A(\ph_segset_h[31] ), 
        .B(seg_cnfg_h) );
    snl_invx05 \BLU/U427  ( .ZN(\BLU/n1548 ), .A(\BLU/n1468 ) );
    snl_invx05 \CODEIF/U266  ( .ZN(\CODEIF/n3875 ), .A(\CODEIF/pfctr[3] ) );
    snl_aoi012x1 \ALUIS/U88  ( .ZN(\ALUIS/n3701 ), .A(\pgldi[5] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_aoi012x1 \LBUS/U560  ( .ZN(\LBUS/*cell*3982/U111/CONTROL2 ), .A(
        \LBUS/MMBSEL ), .B(\LBUS/temp1[2] ), .C(\LBUS/n1399 ) );
    snl_xnor2x0 \CONS/U217  ( .ZN(\CONS/n706 ), .A(\pk_idcz_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_nand13x1 \BLU/U381  ( .ZN(\BLU/n1542 ), .A(\BLU/n1540 ), .B(
        \BLU/n1501 ), .C(\BLU/n1510 ) );
    snl_invx05 \BLU/U400  ( .ZN(\BLU/n1512 ), .A(\pgld16[0] ) );
    snl_muxi21x1 \LDIS/U190  ( .ZN(\LDIS/ldexch[20] ), .A(\LDIS/n3144 ), .B(
        \LDIS/n3143 ), .S(\LDIS/n3165 ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[6]  ( .Q(\pgld32[6] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[6] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_nor02x1 \LBUS/U650  ( .ZN(\LBUS/n1410 ), .A(\LBUS/lnsa_end ), .B(
        \LBUS/n1402 ) );
    snl_and02x1 \REG_2/U146  ( .Z(\ph_cpudout[16] ), .A(\ph_segset_h[16] ), 
        .B(seg_cnfg_h) );
    snl_nand03x0 \CONS/U127  ( .ZN(\CONS/n664 ), .A(\CONS/n665 ), .B(
        ph_bitsrc_h), .C(\CONS/n666 ) );
    snl_ao022x2 \CMPX/U8  ( .Z(ph_lwdsrc_h), .A(ph_lwdsrch), .B(ph_saexe_sth), 
        .C(po_lwdsrc_h), .D(\CMPX/n1047 ) );
    snl_invx05 \REGF/U754  ( .ZN(\REGF/n8192 ), .A(\pgsdprlh[8] ) );
    snl_ao222x1 \CODEIF/U208  ( .Z(\CODEIF/n3855 ), .A(PA[17]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[14] ), .E(cif_byte), .F(PDLIN[14]
        ) );
    snl_invx05 \CONS/U279  ( .ZN(\CONS/n585 ), .A(\CONS/SACO[0] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[12]  ( .Q(\ph_segset_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[12]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_xor2x0 \CODEIF/U398  ( .Z(\CODEIF/n4036 ), .A(\CODEIF/n4035 ), .B(
        \CODEIF/n3992 ) );
    snl_xnor2x0 \CODEIF/U419  ( .ZN(\CODEIF/n4016 ), .A(CDOUT[9]), .B(CDOUT[8]
        ) );
    snl_xor2x0 \LDCHK/U82  ( .Z(\LDCHK/n3270 ), .A(\LDCHK/n3245 ), .B(
        \LDCHK/n3307 ) );
    snl_invx1 \REG_2/U128  ( .ZN(\REG_2/n435 ), .A(\REG_2/n410 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[21]  ( .Q(\ph_segset_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[21]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_invx05 \REGF/U773  ( .ZN(\REGF/n8178 ), .A(\pgsdprlh[15] ) );
    snl_invx05 \ADOSEL/U53  ( .ZN(\ADOSEL/n4108 ), .A(\pkdptout[6] ) );
    snl_nand02x1 \PDOSEL/U145  ( .ZN(\PDOSEL/n117 ), .A(CDIN[25]), .B(
        \PDOSEL/n119 ) );
    snl_nor03x0 \CONS/U149  ( .ZN(\CONS/n523 ), .A(\CONS/n615 ), .B(
        \CONS/n613 ), .C(\CONS/n614 ) );
    snl_and02x1 \REGF/U831  ( .Z(\REGF/n8152 ), .A(\REGF/n8160 ), .B(
        \REGF/n8162 ) );
    snl_invx05 \ADOSEL/U74  ( .ZN(\ADOSEL/n4122 ), .A(\pkdptout[27] ) );
    snl_nor02x1 \LBUS/U619  ( .ZN(\LBUS/n1435 ), .A(\LBUS/n1444 ), .B(
        \LBUS/ilt[5] ) );
    snl_nand02x1 \PDOSEL/U162  ( .ZN(\PDOSEL/n115 ), .A(CDIN[10]), .B(
        \PDOSEL/n119 ) );
    snl_ffqx1 \REGF/D2_HINT_reg  ( .Q(\REGF/D2_HINT ), .D(HINT), .CP(SCLK) );
    snl_invx05 \CODEIF/U283  ( .ZN(\CODEIF/n3906 ), .A(PDLIN[13]) );
    snl_and02x1 \UPIF/U18  ( .Z(\ph_pdis_h[0] ), .A(\pk_rread_h[63] ), .B(
        \UPIF/n1046 ) );
    snl_invx05 \BLU/U364  ( .ZN(\BLU/n1488 ), .A(\pgld16[8] ) );
    snl_xor2x0 \CODEIF/U313  ( .Z(\CODEIF/n3986 ), .A(CDIN[27]), .B(
        \CODEIF/n3985 ) );
    snl_aoi022x1 \ALUIS/U123  ( .ZN(\ALUIS/n3728 ), .A(\stream4[19] ), .B(
        immbsel), .C(\pk_adb_h[19] ), .D(po_brsel_h) );
    snl_xnor2x0 \LDCHK/U106  ( .ZN(\LDCHK/n3283 ), .A(\pgmuxout[20] ), .B(
        \pgmuxout[22] ) );
    snl_muxi21x1 \LDIS/U175  ( .ZN(\LDIS/ldexcl[12] ), .A(\LDIS/n3157 ), .B(
        \LDIS/n3158 ), .S(\LDIS/n3134 ) );
    snl_invx05 \LBUS/U585  ( .ZN(LASOUT), .A(\LBUS/ilt[2] ) );
    snl_nand02x2 \REGF/U375  ( .ZN(\REGF/n8051 ), .A(\REGF/n8228 ), .B(
        ph_tprsel_h) );
    snl_ao2222x1 \REGF/U543  ( .Z(\REGF/RI_SRDA[14] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[14]), .C(\pgldi[14] ), .D(\REGF/n8210 ), .E(\stream3[14] ), .F(
        \REGF/n8211 ), .G(\pkdptout[14] ), .H(\REGF/n8212 ) );
    snl_and02x1 \REGF/U558  ( .Z(\REGF/RO_LPSAS2156[0] ), .A(ph_sastlth), .B(
        \REGF/RO_EST1[0] ) );
    snl_invx05 \REGF/U668  ( .ZN(\REGF/n8189 ), .A(\pgregadrh[9] ) );
    snl_ao222x1 \CODEIF/U194  ( .Z(\CODEIF/n3765 ), .A(cif_cont), .B(PA[3]), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[0] ), .E(cif_byte), .F(PDLIN[0])
         );
    snl_ffandx1 \LBUS/lnsa_err_reg  ( .Q(\LBUS/lnsa_err ), .A(\LBUS/temp[3] ), 
        .B(\LBUS/*cell*3982/U158/Z_0 ), .CP(SCLK) );
    snl_xor2x0 \CONS/U47  ( .Z(\CONS/n569 ), .A(\pk_saco_lh[21] ), .B(
        \pgsdprlh[21] ) );
    snl_sffqenrnx2 \SAEXE/ph_saexe_sth_reg  ( .Q(ph_saexe_sth), .D(1'b0), .EN(
        1'b1), .RN(n10735), .SD(\pk_rwrit_h[49] ), .SE(
        \SAEXE/*cell*3651/U11/CONTROL1 ), .CP(SCLK) );
    snl_nor02x1 \SAEXE/U122  ( .ZN(\SAEXE/singlen ), .A(\pk_psae_h[6] ), .B(
        \pk_psae_h[7] ) );
    snl_invx05 \LDIS/U152  ( .ZN(\LDIS/n3119 ), .A(\pgld32[19] ) );
    snl_oai012x1 \PDOSEL/U36  ( .ZN(PDH[52]), .A(\PDOSEL/n106 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_mux21x1 \ALUSHT/U21  ( .Z(\pkdptout[2] ), .A(\ALUSHT/pkshtout[2] ), 
        .B(\ALUSHT/pkaluout[2] ), .S(\ALUSHT/n3112 ) );
    snl_and02x2 \UPIF/U6  ( .Z(\ph_pdis_h[9] ), .A(\pk_rread_h[42] ), .B(
        \UPIF/n1046 ) );
    snl_oai013x0 \LBUS/U692  ( .ZN(\LBUS/n1607 ), .A(\LBUS/n1456 ), .B(
        \LBUS/n1593 ), .C(\LBUS/ilt[2] ), .D(\LBUS/n1455 ) );
    snl_xor2x0 \CONS/U60  ( .Z(\CONS/n577 ), .A(\CONS/SACO[19] ), .B(
        \pgsdprlh[23] ) );
    snl_xor2x0 \CODEIF/U334  ( .Z(\CODEIF/n4015 ), .A(\CODEIF/n4016 ), .B(
        \CODEIF/n4017 ) );
    snl_aoi012x1 \ALUIS/U104  ( .ZN(\ALUIS/n3745 ), .A(\pgldi[27] ), .B(
        srcbsel), .C(allfbsel) );
    snl_oa012x1 \SAEXE/U105  ( .Z(phrelbwrh), .A(\SAEXE/n416 ), .B(
        \SAEXE/relbwrh ), .C(ph_saexe_sth) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[31]  ( .Q(\pgld32[31] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[31] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_invx05 \BLU/U343  ( .ZN(\BLU/n1558 ), .A(baccsel) );
    snl_invx05 \LDCHK/U121  ( .ZN(\LDCHK/n3267 ), .A(\pgld32[29] ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[28]  ( .Q(\pgld32[28] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[28] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_oai022x1 \REGF/U654  ( .ZN(\REGF/RI_TBAI[0] ), .A(\REGF/n8225 ), .B(
        \REGF/n8138 ), .C(\REGF/n8226 ), .D(\REGF/n8199 ) );
    snl_invx05 \REGF/U673  ( .ZN(\REGF/n8129 ), .A(PDLIN[7]) );
    snl_nand02x1 \ADOSEL/U110  ( .ZN(\ADOSEL/n4124 ), .A(\pgbluext[27] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U76  ( .ZN(\pgaluinb[28] ), .A(\ALUIS/n3746 ), .B(
        \ALUIS/n3747 ) );
    snl_nand03x0 \BLU/U358  ( .ZN(\BLU/n1544 ), .A(\BLU/n1471 ), .B(
        \BLU/n1474 ), .C(\BLU/n1468 ) );
    snl_aoi0b12x0 \LDCHK/U35  ( .ZN(pgldperrh), .A(\LDCHK/n3236 ), .B(
        \LDCHK/n3237 ), .C(\LDCHK/pchkenh ) );
    snl_invx1 \MAIN/U120  ( .ZN(\MAIN/n3611 ), .A(\MAIN/n3610 ) );
    snl_invx05 \LDIS/U149  ( .ZN(\LDIS/n3122 ), .A(\pgld32[22] ) );
    snl_oai012x1 \LBUS/U689  ( .ZN(\LBUS/n1605 ), .A(LDK), .B(\LBUS/n1423 ), 
        .C(\LBUS/n1461 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[31]  ( .Q(\ph_segset_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[31]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[28]  ( .Q(\ph_segset_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[28]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_invx05 \SAEXE/U139  ( .ZN(\SAEXE/n424 ), .A(\pk_psae_h[2] ) );
    snl_oai222x2 \REGF/U390  ( .ZN(\REGF/RI_SRA12M[25] ), .A(\REGF/n8063 ), 
        .B(\REGF/n8051 ), .C(\REGF/n8227 ), .D(\REGF/n8156 ), .E(\REGF/n8228 ), 
        .F(\REGF/n8155 ) );
    snl_oai222x0 \REGF/U458  ( .ZN(\REGF/RI_EACC[7] ), .A(\REGF/n8127 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8128 ), .E(\REGF/n8129 ), 
        .F(\REGF/n8059 ) );
    snl_and02x1 \REGF/U564  ( .Z(\REGF/RO_LPSAS2156[6] ), .A(
        \REGF/RO_PSASL[8] ), .B(ph_sastlth) );
    snl_oai122x0 \CODEIF/U234  ( .ZN(\CODEIF/pfctr415[13] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3905 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3906 ), .E(
        \CODEIF/n3907 ) );
    snl_muxi21x1 \CODEIF/U298  ( .ZN(\CODEIF/write_prtect336 ), .A(
        \CODEIF/n3928 ), .B(\CODEIF/n3866 ), .S(pr_write_h) );
    snl_xor2x0 \CODEIF/U308  ( .Z(\CODEIF/n3978 ), .A(CDIN[38]), .B(
        \CODEIF/n3977 ) );
    snl_nand02x1 \ALUIS/U51  ( .ZN(\pgaluinb[3] ), .A(\ALUIS/n3696 ), .B(
        \ALUIS/n3697 ) );
    snl_aoi012x1 \ALUIS/U138  ( .ZN(\ALUIS/n3713 ), .A(\pgldi[11] ), .B(
        srcbsel), .C(allfbsel) );
    snl_invx05 \CODEIF/U425  ( .ZN(\CODEIF/n4030 ), .A(cnt_write_h) );
    snl_xnor2x0 \CONS/U245  ( .ZN(\CONS/n522 ), .A(\pk_idcy_h[1] ), .B(
        \pk_indy_h[1] ) );
    snl_oai222x0 \REGF/U581  ( .ZN(\REGF/RI_ACC[20] ), .A(\REGF/n8088 ), .B(
        \REGF/n8215 ), .C(\REGF/n8089 ), .D(\REGF/n8216 ), .E(\REGF/n8090 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U721  ( .ZN(\REGF/n8139 ), .A(\pgldi[3] ) );
    snl_invx05 \REGF/U768  ( .ZN(\REGF/n8205 ), .A(\pgregadrh[1] ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[21]  ( .Q(\pgld32[21] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[21] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_aoi022x1 \LBUS/U602  ( .ZN(\LBUS/n1455 ), .A(\LBUS/ilt[5] ), .B(
        \LBUS/ilt[1] ), .C(\LBUS/n1453 ), .D(\LBUS/n1456 ) );
    snl_xnor2x0 \CONS/U175  ( .ZN(\CONS/n652 ), .A(\pgsdprlh[6] ), .B(
        \pk_saco_lh[6] ) );
    snl_oai122x0 \ADOSEL/U26  ( .ZN(\pgmuxout[15] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4134 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4135 ), .E(
        \ADOSEL/n4136 ) );
    snl_invx05 \ADOSEL/U48  ( .ZN(\ADOSEL/n4113 ), .A(\pkdptout[24] ) );
    snl_nor04x0 \CONS/U152  ( .ZN(\CONS/n526 ), .A(\CONS/n722 ), .B(
        \CONS/n618 ), .C(\CONS/n616 ), .D(\CONS/n617 ) );
    snl_invx05 \PDOSEL/U81  ( .ZN(\PDOSEL/n82 ), .A(CDIN[38]) );
    snl_invx1 \CODEIF/U213  ( .ZN(\CODEIF/n3862 ), .A(\CODEIF/n3860 ) );
    snl_xor2x0 \LDCHK/U99  ( .Z(\LDCHK/n3251 ), .A(\LDCHK/n3311 ), .B(
        \LDCHK/pglpinff[1] ) );
    snl_nor02x1 \LBUS/U625  ( .ZN(\LBUS/n1454 ), .A(\LBUS/n1596 ), .B(
        \LBUS/n1597 ) );
    snl_ao022x1 \REG_2/U133  ( .Z(\ph_cpudout[3] ), .A(\ph_segset_h[3] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[3] ), .D(ret_cont_h) );
    snl_xor2x0 \CODEIF/U383  ( .Z(\CODEIF/n4032 ), .A(\CODEIF/n3974 ), .B(
        \CODEIF/n3978 ) );
    snl_xnor2x0 \CODEIF/U402  ( .ZN(\CODEIF/n3996 ), .A(CDOUT[53]), .B(CDOUT
        [55]) );
    snl_xnor2x0 \CONS/U262  ( .ZN(\CONS/n742 ), .A(\pk_idcw_h[20] ), .B(
        \pk_indw_h[20] ) );
    snl_nor02x1 \PDOSEL/U130  ( .ZN(\PDOSEL/n123 ), .A(\ph_cpudout[13] ), .B(
        \pk_pdo_h[13] ) );
    snl_ao022x1 \REGF/U411  ( .Z(\REGF/RI_PCOH[22] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[22]), .C(\stream4[54] ), .D(\REGF/n8053 ) );
    snl_ao2b2b2x0 \REGF/U436  ( .Z(\REGF/RI_EACC[29] ), .A(\REGF/n8063 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8064 ), .E(PDLIN[29]), .F(
        \ph_pdis_h[1] ) );
    snl_aoi022x1 \ALUIS/U93  ( .ZN(\ALUIS/n3696 ), .A(\stream4[3] ), .B(
        immbsel), .C(\pk_adb_h[3] ), .D(po_brsel_h) );
    snl_oai222x0 \REGF/U488  ( .ZN(\REGF/RI_DPR[5] ), .A(\REGF/n8197 ), .B(
        \REGF/n8160 ), .C(\REGF/n8198 ), .D(\REGF/n8162 ), .E(\REGF/n8135 ), 
        .F(\REGF/n8151 ) );
    snl_oai222x0 \REGF/U628  ( .ZN(\REGF/RI_SPR[1] ), .A(\REGF/n8205 ), .B(
        \REGF/n8220 ), .C(\REGF/n8206 ), .D(\REGF/n8221 ), .E(\REGF/n8147 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U696  ( .ZN(\REGF/n8171 ), .A(\pgregadrh[18] ) );
    snl_invx05 \REGF/U706  ( .ZN(\REGF/n8199 ), .A(\pgregadrh[4] ) );
    snl_nor02x1 \PDOSEL/U117  ( .ZN(\PDOSEL/n118 ), .A(\ph_cpudout[25] ), .B(
        \pk_pdo_h[25] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[4]  ( .Q(\REGF/RO_LLPSAS[6] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[4] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_ffqsnx1 \CODEIF/pgfpoel_reg  ( .Q(CROE), .D(\CODEIF/pgfpoe_in ), .SN(
        \CODEIF/n3861 ), .CP(SCLK) );
    snl_xor2x0 \CODEIF/U366  ( .Z(\CODEIF/n3941 ), .A(CDOUT[18]), .B(
        \CODEIF/n4026 ) );
    snl_nand02x1 \ALUIS/U156  ( .ZN(\ALUIS/n3685 ), .A(\pk_ada_h[27] ), .B(
        po_arsel_h) );
    snl_ao022x1 \BLUOS/U26  ( .Z(\pgbluext[7] ), .A(\pkbludgh[7] ), .B(
        ph_bit_h), .C(\pkdptout[7] ), .D(ph_word16_h) );
    snl_and03x1 \CONS/U32  ( .Z(ph_sacons_h), .A(pk_sasea_h), .B(\CONS/n536 ), 
        .C(\CONS/n537 ) );
    snl_ao022x1 \MAIN/U169  ( .Z(\MAIN/n3634 ), .A(sequencial1), .B(
        \MAIN/ph_rdwr1selh ), .C(sequencial2), .D(\MAIN/ph_rdwr2selh ) );
    snl_ao022x1 \LDIS/U100  ( .Z(\pgldi[1] ), .A(ph_word32_h), .B(\pgld32[1] ), 
        .C(\pgld16[1] ), .D(ph_word16_h) );
    snl_or02x1 \CMPX/U11  ( .Z(ph_lbwrh), .A(phrelbwrh), .B(phlbdir) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[3]  ( .Q(\REG_2/ph_retcnt_h[3] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[3]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_oai112x0 \PDOSEL/U64  ( .ZN(PDLOUT[17]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n103 ), .C(\PDOSEL/n152 ), .D(\PDOSEL/n153 ) );
    snl_oai022x1 \BLU/U311  ( .ZN(\pkbludgh[5] ), .A(\BLU/n1464 ), .B(
        \BLU/n1495 ), .C(\BLU/n1496 ), .D(\BLU/n1497 ) );
    snl_nand02x1 \CODEIF/U341  ( .ZN(\CODEIF/n3889 ), .A(\CODEIF/pgctrinc[7] ), 
        .B(\CODEIF/n3945 ) );
    snl_nand02x2 \ALUIS/U18  ( .ZN(\pgaluina[6] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3664 ) );
    snl_nand02x1 \ALUIS/U171  ( .ZN(\ALUIS/n3671 ), .A(\pk_ada_h[13] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U217  ( .ZN(\LDIS/n3159 ), .A(LIN[11]) );
    snl_nor02x1 \BLU/U336  ( .ZN(\BLU/n1481 ), .A(\BLU/n1530 ), .B(\BLU/n1529 
        ) );
    snl_ao022x1 \LDIS/U127  ( .Z(\pgld16[14] ), .A(ph_selldl), .B(\pgld32[14] 
        ), .C(ph_selldh), .D(\pgld32[30] ) );
    snl_xnor2x0 \CONS/U190  ( .ZN(\CONS/n672 ), .A(\pgsdprlh[16] ), .B(
        \CONS/SACO[12] ) );
    snl_oai012x1 \PDOSEL/U43  ( .ZN(PDH[59]), .A(\PDOSEL/n113 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_ao022x1 \LDIS/U112  ( .Z(\pgldi[7] ), .A(ph_word32_h), .B(\pgld32[7] ), 
        .C(\pgld16[7] ), .D(ph_word16_h) );
    snl_nor04x0 \PDOSEL/U76  ( .ZN(\PDOSEL/n223 ), .A(BE[7]), .B(BE[6]), .C(BE
        [4]), .D(BE[5]) );
    snl_ao022x1 \REGF/U518  ( .Z(\REGF/RI_PCOL[7] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[7]), .C(\stream4[7] ), .D(\REGF/n8209 ) );
    snl_invx05 \REGF/U733  ( .ZN(\REGF/n8073 ), .A(\pgldi[25] ) );
    snl_oai122x0 \ADOSEL/U34  ( .ZN(\pgmuxout[23] ), .A(\ADOSEL/n4111 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4110 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4146 ) );
    snl_nand02x1 \ADOSEL/U98  ( .ZN(\ADOSEL/n4145 ), .A(\pgbluext[6] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \CODEIF/U353  ( .ZN(\CODEIF/n3907 ), .A(\CODEIF/pgctrinc[13] 
        ), .B(\CODEIF/n3945 ) );
    snl_xnor2x0 \CODEIF/U374  ( .ZN(\CODEIF/n3968 ), .A(CDIN[52]), .B(CPIN[3])
         );
    snl_nand02x1 \ALUIS/U144  ( .ZN(\ALUIS/n3667 ), .A(po_arsel_h), .B(
        \pk_ada_h[9] ) );
    snl_oai022x1 \BLU/U303  ( .ZN(\pkbludgh[13] ), .A(\BLU/n1464 ), .B(
        \BLU/n1471 ), .C(\BLU/n1472 ), .D(\BLU/n1473 ) );
    snl_nand02x1 \ALUIS/U163  ( .ZN(\ALUIS/n3678 ), .A(\pk_ada_h[20] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U222  ( .ZN(\LDIS/n3156 ), .A(LIN[29]) );
    snl_sffqrnx1 \LBUS/flag_tr2_reg  ( .Q(\LBUS/flag_tr2 ), .D(1'b0), .RN(
        n10734), .SD(\LBUS/n1393 ), .SE(pgoddflgh), .CP(SCLK) );
    snl_ao022x1 \BLUOS/U13  ( .Z(\pgbluext[16] ), .A(\pkbludgh[0] ), .B(
        ph_bit_h), .C(\pkdptout[0] ), .D(ph_word16_h) );
    snl_aoi022x1 \LDCHK/U49  ( .ZN(\LDCHK/n3266 ), .A(\LDCHK/n3267 ), .B(
        \LDCHK/n3255 ), .C(\pgld32[29] ), .D(\pgld32[31] ) );
    snl_invx05 \LDIS/U205  ( .ZN(\LDIS/n3141 ), .A(LIN[5]) );
    snl_nor02x1 \BLU/U324  ( .ZN(\BLU/n1490 ), .A(\BLU/n1533 ), .B(\BLU/n1534 
        ) );
    snl_ao022x1 \CMPX/U24  ( .Z(ph_sais_h), .A(\CMPX/n1051 ), .B(ph_saexe_sth), 
        .C(po_trsset_h), .D(\CMPX/n1047 ) );
    snl_oai012x1 \LDIS/U135  ( .ZN(\pgldi[21] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3121 ), .C(\LDIS/n3115 ) );
    snl_invx05 \LDIS/U199  ( .ZN(\LDIS/n3147 ), .A(LIN[2]) );
    snl_xnor2x0 \CONS/U182  ( .ZN(\CONS/n659 ), .A(\pgsdprlh[16] ), .B(
        \pk_saco_lh[16] ) );
    snl_ao112x1 \PDOSEL/U51  ( .Z(PDLOUT[28]), .A(CDIN[28]), .B(\PDOSEL/n119 ), 
        .C(\pk_pdo_h[28] ), .D(\ph_cpudout[28] ) );
    snl_nor02x1 \PDOSEL/U122  ( .ZN(\PDOSEL/n125 ), .A(\ph_cpudout[20] ), .B(
        \pk_pdo_h[20] ) );
    snl_nand03x0 \LBUS/U659  ( .ZN(\LBUS/n1414 ), .A(
        \LBUS/*cell*3982/U71/CONTROL1 ), .B(\LBUS/n1439 ), .C(stage_a) );
    snl_nand02x1 \BLU/U388  ( .ZN(\BLU/n1465 ), .A(\BLU/n1567 ), .B(
        \BLU/n1565 ) );
    snl_and02x1 \BLU/U409  ( .Z(\BLU/n1582 ), .A(pkalucmf), .B(\BLU/n1558 ) );
    snl_oai2222x0 \REGF/U367  ( .ZN(\REGF/RI_SRA12M[2] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8144 ), .C(\REGF/n8142 ), .D(\REGF/n8051 ), .E(\REGF/n8229 ), 
        .F(\REGF/n8203 ), .G(\REGF/n8230 ), .H(\REGF/n8204 ) );
    snl_oai2222x0 \REGF/U382  ( .ZN(\REGF/RI_SRA12M[4] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8138 ), .C(\REGF/n8136 ), .D(\REGF/n8051 ), .E(\REGF/n8199 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8200 ) );
    snl_invx1 \REGF/U403  ( .ZN(\REGF/n8151 ), .A(\ph_pdis_h[2] ) );
    snl_ao022x1 \REGF/U424  ( .Z(\REGF/RI_PCOH[9] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[9]), .C(\REGF/n8053 ), .D(\stream4[41] ) );
    snl_oai222x0 \REGF/U593  ( .ZN(\REGF/RI_ACC[8] ), .A(\REGF/n8124 ), .B(
        \REGF/n8215 ), .C(\REGF/n8125 ), .D(\REGF/n8216 ), .E(\REGF/n8126 ), 
        .F(\REGF/n8217 ) );
    snl_xor2x0 \CODEIF/U248  ( .Z(CPOUT[0]), .A(\CODEIF/n3942 ), .B(
        \CODEIF/n3943 ) );
    snl_aoi022x1 \ALUIS/U81  ( .ZN(\ALUIS/n3708 ), .A(immbsel), .B(
        \stream4[9] ), .C(po_brsel_h), .D(\pk_adb_h[9] ) );
    snl_nand02x1 \LBUS/U569  ( .ZN(\LBUS/*cell*3982/U200/CONTROL1 ), .A(
        \LBUS/n1400 ), .B(\LBUS/n1414 ) );
    snl_xnor2x0 \CONS/U239  ( .ZN(\CONS/n725 ), .A(\pk_idcy_h[20] ), .B(
        \pk_indy_h[20] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[16]  ( .Q(\ph_segset_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[16]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_ao2222x1 \REGF/U551  ( .Z(\REGF/RI_SRDA[6] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[6]), .C(\pgldi[6] ), .D(\REGF/n8210 ), .E(\stream3[6] ), .F(
        \REGF/n8211 ), .G(\pkdptout[6] ), .H(\REGF/n8212 ) );
    snl_invx05 \REGF/U684  ( .ZN(\REGF/n8197 ), .A(\pgregadrh[5] ) );
    snl_oai122x0 \ADOSEL/U13  ( .ZN(\pgmuxout[2] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4095 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4096 ), .E(
        \ADOSEL/n4097 ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[12]  ( .Q(\pgld32[12] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexcl[12] ), .SE(lo_data_lth), .CP(SCLK
        ) );
    snl_xor2x0 \CONS/U109  ( .Z(\CONS/n627 ), .A(\pk_idcx_h[15] ), .B(
        \pk_indx_h[15] ) );
    snl_invx05 \PDOSEL/U105  ( .ZN(\PDOSEL/n74 ), .A(CDIN[32]) );
    snl_invx05 \REGF/U714  ( .ZN(\REGF/n8121 ), .A(\pgldi[9] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[9]  ( .Q(\REGF/RO_LLPSAS[13] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[9] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_ao222x1 \CODEIF/U201  ( .Z(\CODEIF/n3848 ), .A(PA[10]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[7] ), .E(cif_byte), .F(PDLIN[7])
         );
    snl_oai122x0 \CODEIF/U226  ( .ZN(\CODEIF/pfctr415[5] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3881 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3882 ), .E(
        \CODEIF/n3883 ) );
    snl_xnor2x0 \CONS/U257  ( .ZN(\CONS/n351 ), .A(\pk_idcx_h[10] ), .B(
        \pk_indx_h[10] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[25]  ( .Q(\ph_segset_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[25]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_muxi21x1 \BLU/U440  ( .ZN(\BLU/n1587 ), .A(\BLU/n1577 ), .B(
        \BLU/n1578 ), .S(\poalufnc[3] ) );
    snl_xnor2x0 \CODEIF/U391  ( .ZN(\CODEIF/n4034 ), .A(CDIN[15]), .B(CDIN[18]
        ) );
    snl_xor2x0 \CODEIF/U410  ( .Z(\CODEIF/n4025 ), .A(\CODEIF/n4039 ), .B(
        CDOUT[39]) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[2]  ( .Q(\pgld32[2] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[2] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_nand12x1 \CONS/U167  ( .ZN(\CONS/n536 ), .A(ph_atchkenh), .B(
        pk_sased_h) );
    snl_nor02x1 \LBUS/U610  ( .ZN(\LBUS/n1460 ), .A(\LBUS/ilt[4] ), .B(
        \LBUS/ilt[5] ) );
    snl_invx05 \LBUS/U637  ( .ZN(\LBUS/n1458 ), .A(LBER) );
    snl_nand02x1 \CONS/U140  ( .ZN(\CONS/n699 ), .A(\CONS/n700 ), .B(
        \CONS/n701 ) );
    snl_invx05 \PDOSEL/U93  ( .ZN(\PDOSEL/n106 ), .A(CDIN[52]) );
    snl_xnor2x0 \CONS/U270  ( .ZN(\CONS/n342 ), .A(\pk_idcw_h[13] ), .B(
        \pk_indw_h[13] ) );
    snl_oai222x0 \REGF/U576  ( .ZN(\REGF/RI_ACC[25] ), .A(\REGF/n8073 ), .B(
        \REGF/n8215 ), .C(\REGF/n8074 ), .D(\REGF/n8216 ), .E(\REGF/n8075 ), 
        .F(\REGF/n8217 ) );
    snl_oai022x1 \REGF/U646  ( .ZN(\REGF/RI_TBAI[8] ), .A(\REGF/n8225 ), .B(
        \REGF/n8114 ), .C(\REGF/n8226 ), .D(\REGF/n8183 ) );
    snl_invx05 \REGF/U661  ( .ZN(\REGF/n8111 ), .A(PDLIN[13]) );
    snl_nand02x1 \ADOSEL/U102  ( .ZN(\ADOSEL/n4142 ), .A(\pgbluext[3] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U64  ( .ZN(\pgaluinb[16] ), .A(\ALUIS/n3722 ), .B(
        \ALUIS/n3723 ) );
    snl_mux21x1 \ALUSHT/U28  ( .Z(\pkdptout[23] ), .A(\ALUSHT/pkshtout[23] ), 
        .B(\ALUSHT/pkaluout[23] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U69  ( .Z(\CONS/n587 ), .A(\pk_pc_h[3] ), .B(
        \pk_pcs2_h[3] ) );
    snl_nand12x1 \MAIN/U132  ( .ZN(\MAIN/ADROVH ), .A(\MAIN/LBAOVFH ), .B(
        \MAIN/n3626 ) );
    snl_oai012x1 \PDOSEL/U18  ( .ZN(PDH[34]), .A(\PDOSEL/n78 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_oai222x0 \REGF/U476  ( .ZN(\REGF/RI_DPR[17] ), .A(\REGF/n8173 ), .B(
        \REGF/n8160 ), .C(\REGF/n8174 ), .D(\REGF/n8162 ), .E(\REGF/n8099 ), 
        .F(\REGF/n8151 ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[0]  ( .Q(\REGF/RO_LLPSAS[0] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[0] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_nand02x1 \ALUIS/U43  ( .ZN(\pgaluina[27] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3685 ) );
    snl_and02x1 \UPIF/U11  ( .Z(\ph_pdis_h[3] ), .A(\pk_rread_h[60] ), .B(
        \UPIF/n1046 ) );
    snl_xor2x0 \CODEIF/U291  ( .Z(\CODEIF/n3946 ), .A(\CODEIF/n3947 ), .B(
        \CODEIF/n3948 ) );
    snl_xor2x0 \CODEIF/U301  ( .Z(\CODEIF/n3966 ), .A(\CODEIF/n3967 ), .B(
        \CODEIF/n3968 ) );
    snl_aoi022x1 \ALUIS/U131  ( .ZN(\ALUIS/n3720 ), .A(\stream4[15] ), .B(
        immbsel), .C(\pk_adb_h[15] ), .D(po_brsel_h) );
    snl_nand02x1 \ALUIS/U58  ( .ZN(\pgaluinb[10] ), .A(\ALUIS/n3710 ), .B(
        \ALUIS/n3711 ) );
    snl_invx05 \BLU/U376  ( .ZN(\BLU/n1500 ), .A(\pgld16[4] ) );
    snl_xor2x0 \CODEIF/U326  ( .Z(\CODEIF/n4005 ), .A(CDOUT[36]), .B(
        \CODEIF/n4004 ) );
    snl_aoi012x1 \ALUIS/U116  ( .ZN(\ALUIS/n3733 ), .A(\pgldi[21] ), .B(
        srcbsel), .C(allfbsel) );
    snl_aoi013x0 \MAIN/U129  ( .ZN(\MAIN/seq_enable ), .A(\MAIN/n3620 ), .B(
        \MAIN/n3621 ), .C(\MAIN/n3622 ), .D(\MAIN/n3623 ) );
    snl_xnor2x0 \LDCHK/U114  ( .ZN(\LDCHK/n3291 ), .A(\pgmuxout[7] ), .B(
        \pgmuxout[5] ) );
    snl_nor02x1 \LBUS/U597  ( .ZN(\LBUS/n1450 ), .A(LDK), .B(\LBUS/n1423 ) );
    snl_oai012x1 \LDIS/U140  ( .ZN(\pgldi[26] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3126 ), .C(\LDIS/n3115 ) );
    snl_muxi21x1 \LDIS/U167  ( .ZN(\LDIS/ldexcl[5] ), .A(\LDIS/n3141 ), .B(
        \LDIS/n3142 ), .S(\LDIS/n3134 ) );
    snl_ffqrnx1 \LBUS/ilt_reg[3]  ( .Q(\LBUS/temp[3] ), .D(\LBUS/nlt[3] ), 
        .RN(n10734), .CP(SCLK) );
    snl_mux21x1 \ALUSHT/U14  ( .Z(\pkdptout[7] ), .A(\ALUSHT/pkshtout[7] ), 
        .B(\ALUSHT/pkaluout[7] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U55  ( .Z(\CONS/n565 ), .A(\CONS/SACO[1] ), .B(
        \pgsdprlh[5] ) );
    snl_invx05 \SAEXE/U130  ( .ZN(\SAEXE/n425 ), .A(\SAEXE/rf_srcadr2_h ) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[7]  ( .Q(\REG_2/ph_retcnt_h[7] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[7]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_oai012x1 \PDOSEL/U24  ( .ZN(PDH[40]), .A(\PDOSEL/n94 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_mux21x1 \ALUSHT/U33  ( .Z(\pkdptout[19] ), .A(\ALUSHT/pkshtout[19] ), 
        .B(\ALUSHT/pkaluout[19] ), .S(\ALUSHT/n3112 ) );
    snl_invx05 \LBUS/U680  ( .ZN(\LBUS/n1609 ), .A(\LBUS/n1457 ) );
    snl_or02x1 \SAEXE/U117  ( .Z(\SAEXE/seq_end ), .A(\SAEXE/exec_end2 ), .B(
        \SAEXE/exec_end1 ) );
    snl_xor2x0 \CONS/U72  ( .Z(\CONS/n590 ), .A(\pk_pcs2_h[12] ), .B(
        \pk_pc_h[12] ) );
    snl_invx05 \BLU/U351  ( .ZN(\BLU/n1566 ), .A(\pgbitnoh[2] ) );
    snl_invx05 \REGF/U804  ( .ZN(\REGF/n8092 ), .A(\pkdptout[19] ) );
    snl_invx1 U10 ( .ZN(n10735), .A(n10737) );
    snl_nand02x2 \REGF/U399  ( .ZN(\REGF/n8221 ), .A(po_ptrsel_h), .B(
        \REGF/n8218 ) );
    snl_oai222x0 \REGF/U451  ( .ZN(\REGF/RI_EACC[14] ), .A(\REGF/n8106 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8107 ), .E(\REGF/n8108 ), 
        .F(\REGF/n8059 ) );
    snl_invx05 \REGF/U746  ( .ZN(\REGF/n8103 ), .A(\pgldi[15] ) );
    snl_invx05 \REGF/U761  ( .ZN(\REGF/n8204 ), .A(\pgsdprlh[2] ) );
    snl_oai122x0 \ADOSEL/U41  ( .ZN(\pgmuxout[30] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4132 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4131 ), .E(
        \ADOSEL/n4153 ) );
    snl_invx05 \LDCHK/U90  ( .ZN(\LDCHK/n3275 ), .A(LPIN[2]) );
    snl_invx05 \PDOSEL/U88  ( .ZN(\PDOSEL/n111 ), .A(CDIN[57]) );
    snl_nand02x1 \PDOSEL/U157  ( .ZN(\PDOSEL/n182 ), .A(CDIN[15]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \ADOSEL/U66  ( .ZN(\ADOSEL/n4131 ), .A(\pkdptout[30] ) );
    snl_nand04x0 \REGF/U823  ( .ZN(\REGF/n8236 ), .A(\REGF/RO_ACC[23] ), .B(
        \REGF/RO_ACC[22] ), .C(\REGF/RO_ACC[20] ), .D(\REGF/RO_ACC[27] ) );
    snl_invx05 \CODEIF/U253  ( .ZN(\CODEIF/n3893 ), .A(\CODEIF/pfctr[9] ) );
    snl_ffqrnx1 \CODEIF/write_prtect_reg  ( .Q(\CODEIF/write_prtect ), .D(
        \CODEIF/write_prtect336 ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_mux21x2 \SHTCD/U10  ( .Z(\phshtd[0] ), .A(\pgld16[0] ), .B(
        \stream4[0] ), .S(immbsel) );
    snl_nor02x2 \LBUS/U555  ( .ZN(lo_data_lth), .A(\LBUS/n1412 ), .B(
        \LBUS/n1437 ) );
    snl_nor03x0 \LBUS/U665  ( .ZN(\LBUS/*cell*3982/U188/CONTROL1 ), .A(
        \LBUS/n1457 ), .B(ph_lbwrh), .C(\LBUS/n1430 ) );
    snl_xor2x0 \CONS/U97  ( .Z(\CONS/n615 ), .A(\pk_idcy_h[11] ), .B(
        \pk_indy_h[11] ) );
    snl_xor2x0 \CONS/U112  ( .Z(\CONS/n630 ), .A(\pk_idcw_h[0] ), .B(
        \pk_indw_h[0] ) );
    snl_oai133x0 \LBUS/U572  ( .ZN(\LBUS/nlt[0] ), .A(\LBUS/n1423 ), .B(
        \LBUS/n1424 ), .C(\LBUS/n1425 ), .D(\LBUS/n1419 ), .E(\LBUS/ilt[0] ), 
        .F(\LBUS/ilt[4] ), .G(\LBUS/n1426 ) );
    snl_xnor2x0 \CONS/U222  ( .ZN(\CONS/n712 ), .A(\pk_idcz_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_invx05 \BLU/U435  ( .ZN(\BLU/n1552 ), .A(\BLU/n1524 ) );
    snl_ao022x1 \REGF/U418  ( .Z(\REGF/RI_PCOH[15] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[15]), .C(\stream4[47] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U438  ( .ZN(\REGF/RI_EACC[27] ), .A(\REGF/n8067 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8068 ), .E(\REGF/n8069 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U493  ( .ZN(\REGF/RI_DPR[0] ), .A(\REGF/n8207 ), .B(
        \REGF/n8160 ), .C(\REGF/n8208 ), .D(\REGF/n8162 ), .E(\REGF/n8150 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U524  ( .Z(\REGF/RI_PCOL[1] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[1]), .C(\stream4[1] ), .D(\REGF/n8209 ) );
    snl_oai222x0 \REGF/U588  ( .ZN(\REGF/RI_ACC[13] ), .A(\REGF/n8109 ), .B(
        \REGF/n8215 ), .C(\REGF/n8110 ), .D(\REGF/n8216 ), .E(\REGF/n8111 ), 
        .F(\REGF/n8217 ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[25]  ( .Q(\pgld32[25] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[25] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_oai222x0 \REGF/U614  ( .ZN(\REGF/RI_SPR[15] ), .A(\REGF/n8177 ), .B(
        \REGF/n8220 ), .C(\REGF/n8178 ), .D(\REGF/n8221 ), .E(\REGF/n8105 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U728  ( .ZN(\REGF/n8065 ), .A(\pgldi[28] ) );
    snl_invx05 \CODEIF/U274  ( .ZN(\CODEIF/n3917 ), .A(\CODEIF/pfctr[17] ) );
    snl_and02x1 \REG_2/U154  ( .Z(\ph_cpudout[24] ), .A(\ph_segset_h[24] ), 
        .B(seg_cnfg_h) );
    snl_nand02x1 \BLU/U393  ( .ZN(\BLU/n1471 ), .A(\BLU/n1570 ), .B(
        \BLU/n1567 ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[16]  ( .Q(\pgld32[16] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[16] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_xnor2x0 \CONS/U205  ( .ZN(\CONS/n688 ), .A(\pk_pc_h[5] ), .B(
        \pk_pcs2_h[5] ) );
    snl_nor03x0 \BLU/U412  ( .ZN(\BLU/n1586 ), .A(allfasel), .B(all0asel), .C(
        all0bsel) );
    snl_nand02x1 \ADOSEL/U83  ( .ZN(\ADOSEL/n4112 ), .A(\pgbluext[7] ), .B(
        \ADOSEL/n4156 ) );
    snl_aoi022x1 \MAIN/U147  ( .ZN(\MAIN/n3631 ), .A(ronly1), .B(
        \MAIN/ph_rdwr1selh ), .C(ronly2), .D(\MAIN/ph_rdwr2selh ) );
    snl_muxi21x1 \LDIS/U182  ( .ZN(\LDIS/ldexch[28] ), .A(\LDIS/n3158 ), .B(
        \LDIS/n3157 ), .S(\LDIS/n3165 ) );
    snl_invx05 \LBUS/U642  ( .ZN(\LBUS/n1419 ), .A(ph_lbussth) );
    snl_nand02x1 \PDOSEL/U139  ( .ZN(\PDOSEL/n162 ), .A(CDIN[5]), .B(
        \PDOSEL/n119 ) );
    snl_nand03x0 \CONS/U135  ( .ZN(\CONS/n682 ), .A(\CONS/n683 ), .B(
        \CONS/n684 ), .C(\CONS/n685 ) );
    snl_xnor2x0 \CONS/U199  ( .ZN(\CONS/n678 ), .A(\pk_pc_h[16] ), .B(
        \pk_pcs2_h[16] ) );
    snl_muxi21x1 \LDCHK/U52  ( .ZN(\LDCHK/lpex[3] ), .A(\LDCHK/n3272 ), .B(
        \LDCHK/n3273 ), .S(\LDCHK/n3274 ) );
    snl_invx05 \REGF/U784  ( .ZN(\REGF/n8125 ), .A(\pkdptout[8] ) );
    snl_nand02x1 \CODEIF/U348  ( .ZN(\CODEIF/n3922 ), .A(\CODEIF/pgctrinc[18] 
        ), .B(\CODEIF/n3945 ) );
    snl_invx1 \ALUIS/U11  ( .ZN(\pgaluina[2] ), .A(\ALUIS/n3643 ) );
    snl_nand02x1 \ALUIS/U36  ( .ZN(\pgaluina[20] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3678 ) );
    snl_nand12x1 \BLU/U318  ( .ZN(ociff), .A(\BLU/n1517 ), .B(\BLU/n1518 ) );
    snl_ao022x1 \REGF/U503  ( .Z(\REGF/RI_PCOL[22] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[22]), .C(\stream4[22] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U633  ( .Z(\REGF/RI_STAT[2] ), .A(\ph_pdis_h[4] ), .B(
        PDLIN[16]), .C(ociff), .D(\REGF/n8224 ) );
    snl_nand02x1 \MAIN/U160  ( .ZN(\MAIN/n3614 ), .A(ciffsel), .B(ph_filewr_h)
         );
    snl_ao022x1 \LDIS/U109  ( .Z(\pgld16[5] ), .A(ph_selldl), .B(\pgld32[5] ), 
        .C(ph_selldh), .D(\pgld32[21] ) );
    snl_invx05 \CMPX/U18  ( .ZN(\CMPX/n1047 ), .A(ph_saexe_sth) );
    snl_oai122x0 \ADOSEL/U28  ( .ZN(\pgmuxout[17] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4093 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4092 ), .E(
        \ADOSEL/n4140 ) );
    snl_xor2x0 \LDCHK/U75  ( .Z(\LDCHK/n3303 ), .A(\pgld32[18] ), .B(
        \pgld32[23] ) );
    snl_or08x1 \CONS/U132  ( .Z(\CONS/n567 ), .A(\CONS/n580 ), .B(\CONS/n581 ), 
        .C(\CONS/n582 ), .D(\CONS/n583 ), .E(\CONS/n584 ), .F(\CONS/n578 ), 
        .G(\CONS/n579 ), .H(\CONS/n552 ) );
    snl_invx05 \CODEIF/U254  ( .ZN(\CODEIF/n3894 ), .A(PDLIN[9]) );
    snl_invx05 \CODEIF/U273  ( .ZN(\CODEIF/n3921 ), .A(PDLIN[18]) );
    snl_muxi21x1 \LDIS/U185  ( .ZN(\LDIS/ldexch[25] ), .A(\LDIS/n3133 ), .B(
        \LDIS/n3132 ), .S(\LDIS/n3165 ) );
    snl_oai012x1 \LBUS/U645  ( .ZN(\LBUS/n1401 ), .A(\LBUS/flag_tr2 ), .B(
        pgoddflgh), .C(ph_lbussth) );
    snl_and02x1 \REG_2/U153  ( .Z(\ph_cpudout[23] ), .A(\ph_segset_h[23] ), 
        .B(seg_cnfg_h) );
    snl_nand04x0 \LBUS/U575  ( .ZN(\LBUS/nlt[4] ), .A(\LBUS/n1397 ), .B(
        \LBUS/n1431 ), .C(\LBUS/n1432 ), .D(\LBUS/n1433 ) );
    snl_xnor2x0 \CONS/U202  ( .ZN(\CONS/n685 ), .A(\pk_pc_h[9] ), .B(
        \pk_pcs2_h[9] ) );
    snl_oa2222x1 \BLU/U415  ( .Z(\BLU/n1514 ), .A(\BLU/n1486 ), .B(\BLU/n1488 
        ), .C(\BLU/n1483 ), .D(\BLU/n1485 ), .E(\BLU/n1480 ), .F(\BLU/n1482 ), 
        .G(\BLU/n1477 ), .H(\BLU/n1479 ) );
    snl_invx05 \BLU/U394  ( .ZN(\BLU/n1476 ), .A(\pgld16[12] ) );
    snl_sffqenrnx1 \LBUS/EXTSEL_reg  ( .Q(\LBUS/EXTSEL ), .D(1'b0), .EN(1'b1), 
        .RN(n10734), .SD(ph_extselh), .SE(\LBUS/n1393 ), .CP(SCLK) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[27]  ( .Q(\pgld32[27] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[27] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_xnor2x0 \CONS/U225  ( .ZN(\CONS/n532 ), .A(\pk_idcz_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \BLU/U432  ( .ZN(\BLU/n1526 ), .A(allfasel) );
    snl_oai222x0 \REGF/U456  ( .ZN(\REGF/RI_EACC[9] ), .A(\REGF/n8121 ), .B(
        \REGF/n8055 ), .C(\REGF/n8122 ), .D(\REGF/n8056 ), .E(\REGF/n8123 ), 
        .F(\REGF/n8059 ) );
    snl_ao022x1 \REGF/U494  ( .Z(\REGF/RI_PCOL[31] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[31]), .C(\stream4[31] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U504  ( .Z(\REGF/RI_PCOL[21] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[21]), .C(\stream4[21] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U634  ( .Z(\REGF/RI_STAT[1] ), .A(PDLIN[1]), .B(
        \ph_pdis_h[4] ), .C(oebacc), .D(\REGF/n8224 ) );
    snl_invx05 \REGF/U698  ( .ZN(\REGF/n8173 ), .A(\pgregadrh[17] ) );
    snl_nand02x1 \REGF/U708  ( .ZN(\REGF/n8232 ), .A(ph_rgfile_h), .B(
        \REGF/n8223 ) );
    snl_invx1 \LBUS/U552  ( .ZN(ad_latch), .A(\LBUS/n1392 ) );
    snl_nor02x1 \LBUS/U662  ( .ZN(\LBUS/*cell*3982/U119/CONTROL1 ), .A(
        \LBUS/n1401 ), .B(\LBUS/n1439 ) );
    snl_xor2x0 \CONS/U115  ( .Z(\CONS/n633 ), .A(\pk_idcw_h[3] ), .B(
        \pk_indw_h[3] ) );
    snl_nor02x1 \PDOSEL/U119  ( .ZN(\PDOSEL/n177 ), .A(\ph_cpudout[23] ), .B(
        \pk_pdo_h[23] ) );
    snl_xor2x0 \CONS/U90  ( .Z(\CONS/n608 ), .A(\pk_idcz_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_ao022x1 \BLUOS/U28  ( .Z(\pgbluext[9] ), .A(ph_bit_h), .B(
        \pkbludgh[9] ), .C(ph_word16_h), .D(\pkdptout[9] ) );
    snl_xor2x0 \LDCHK/U72  ( .Z(\LDCHK/n3301 ), .A(\pgld32[19] ), .B(
        \pgld32[20] ) );
    snl_invx05 \MAIN/U167  ( .ZN(ph_rmw2h), .A(\MAIN/n3621 ) );
    snl_ao022x1 \REGF/U523  ( .Z(\REGF/RI_PCOL[2] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[2]), .C(\stream4[2] ), .D(\REGF/n8209 ) );
    snl_xor2x0 \CODEIF/U368  ( .Z(\CODEIF/n3943 ), .A(CDOUT[5]), .B(
        \CODEIF/n4028 ) );
    snl_nand02x1 \ALUIS/U31  ( .ZN(\ALUIS/n3754 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3661 ) );
    snl_nand02x1 \ALUIS/U158  ( .ZN(\ALUIS/n3683 ), .A(\pk_ada_h[25] ), .B(
        po_arsel_h) );
    snl_oai222x0 \REGF/U613  ( .ZN(\REGF/RI_SPR[16] ), .A(\REGF/n8175 ), .B(
        \REGF/n8220 ), .C(\REGF/n8176 ), .D(\REGF/n8221 ), .E(\REGF/n8102 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U783  ( .ZN(\REGF/n8122 ), .A(\pkdptout[9] ) );
    snl_and02x1 \ALUIS/U16  ( .Z(\ALUIS/n3649 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3672 ) );
    snl_aoi022x1 \BLU/U338  ( .ZN(\BLU/n1522 ), .A(\BLU/n1552 ), .B(
        \BLU/n1525 ), .C(\BLU/n1524 ), .D(\BLU/n1519 ) );
    snl_muxi21x1 \LDCHK/U55  ( .ZN(\LDCHK/lpex[0] ), .A(\LDCHK/n3276 ), .B(
        \LDCHK/n3275 ), .S(\LDCHK/n3277 ) );
    snl_invx05 \LDIS/U219  ( .ZN(\LDIS/n3157 ), .A(LIN[12]) );
    snl_nand04x0 \REGF/U824  ( .ZN(\REGF/n8237 ), .A(\REGF/RO_ACC[16] ), .B(
        \REGF/RO_ACC[24] ), .C(\REGF/RO_ACC[21] ), .D(\REGF/RO_ACC[18] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[2]  ( .Q(\REGF/RO_LLPSAS[4] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[2] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_nand02x1 \ADOSEL/U84  ( .ZN(\ADOSEL/n4109 ), .A(\pgbluext[6] ), .B(
        \ADOSEL/n4156 ) );
    snl_ao022x1 \LDIS/U129  ( .Z(\pgld16[15] ), .A(ph_selldl), .B(\pgld32[15] 
        ), .C(ph_selldh), .D(\pgld32[31] ) );
    snl_xor2x0 \CODEIF/U321  ( .Z(\CODEIF/n3998 ), .A(CDOUT[50]), .B(
        \CODEIF/n3997 ) );
    snl_nand02x1 \ALUIS/U78  ( .ZN(\pgaluinb[30] ), .A(\ALUIS/n3750 ), .B(
        \ALUIS/n3751 ) );
    snl_aoi022x1 \MAIN/U140  ( .ZN(\MAIN/n3620 ), .A(rmw11), .B(
        \MAIN/ph_rdwr1selh ), .C(rmw12), .D(\MAIN/ph_rdwr2selh ) );
    snl_ffqrnx1 \MAIN/cstregw_tap2_reg  ( .Q(\MAIN/cstregw_tap2 ), .D(
        \MAIN/cstregw_tap1 ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_aoi022x1 \ALUIS/U111  ( .ZN(\ALUIS/n3738 ), .A(\stream4[24] ), .B(
        immbsel), .C(\pk_adb_h[24] ), .D(po_brsel_h) );
    snl_nand03x0 \BLU/U356  ( .ZN(\BLU/n1539 ), .A(\BLU/n1507 ), .B(
        \BLU/n1510 ), .C(\BLU/n1504 ) );
    snl_xor2x0 \CODEIF/U296  ( .Z(\CODEIF/n3959 ), .A(\CODEIF/n3960 ), .B(CPIN
        [0]) );
    snl_xnor2x0 \LDCHK/U113  ( .ZN(\LDCHK/n3290 ), .A(\pgmuxout[3] ), .B(
        \pgmuxout[6] ) );
    snl_invx05 \LDIS/U147  ( .ZN(\LDIS/n3124 ), .A(\pgld32[24] ) );
    snl_mux21x1 \ALUSHT/U34  ( .Z(\pkdptout[18] ), .A(\ALUSHT/pkshtout[18] ), 
        .B(\ALUSHT/pkaluout[18] ), .S(\ALUSHT/n3112 ) );
    snl_invx05 \LBUS/U687  ( .ZN(\LBUS/n1405 ), .A(ph_lbend) );
    snl_xor2x0 \CONS/U75  ( .Z(\CONS/n593 ), .A(\pk_pc_h[13] ), .B(
        \pk_pcs1_h[13] ) );
    snl_oai012x1 \PDOSEL/U23  ( .ZN(PDH[39]), .A(\PDOSEL/n92 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nor02x1 \SAEXE/U110  ( .ZN(ph_srcsl_h), .A(\SAEXE/srcwrit ), .B(
        \SAEXE/n413 ) );
    snl_invx05 \LDIS/U160  ( .ZN(\LDIS/n3126 ), .A(\pgld32[26] ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[9]  ( .Q(\pgld32[9] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[9] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_ffqrnx1 \LBUS/ilt_reg[1]  ( .Q(\LBUS/ilt[1] ), .D(\LBUS/nlt[1] ), .RN(
        n10734), .CP(SCLK) );
    snl_mux21x1 \ALUSHT/U13  ( .Z(\pkdptout[8] ), .A(\ALUSHT/pkshtout[8] ), 
        .B(\ALUSHT/pkaluout[8] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U52  ( .Z(\CONS/n574 ), .A(\pk_saco_lh[1] ), .B(
        \pgsdprlh[1] ) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[5]  ( .Q(\REG_2/ph_retcnt_h[5] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[5]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_invx05 \SAEXE/U137  ( .ZN(\SAEXE/n422 ), .A(\pk_psae_h[4] ) );
    snl_nor04x0 \LBUS/U590  ( .ZN(ph_wdstenh), .A(ph_wdsrdaselh), .B(LRQ), .C(
        \LBUS/n1447 ), .D(\LBUS/n1441 ) );
    snl_sffqenrnx1 \LBUS/word32odphase_reg  ( .Q(\LBUS/word32odphase ), .D(
        1'b0), .EN(1'b1), .RN(n10734), .SD(\LBUS/*cell*3982/U71/CONTROL1 ), 
        .SE(\LBUS/*cell*3982/U176/CONTROL1 ), .CP(SCLK) );
    snl_xor2x0 \CODEIF/U306  ( .Z(\CODEIF/n3974 ), .A(\CODEIF/n3975 ), .B(
        \CODEIF/n3976 ) );
    snl_nand13x1 \BLU/U371  ( .ZN(\BLU/n1536 ), .A(\BLU/n1534 ), .B(
        \BLU/n1489 ), .C(\BLU/n1498 ) );
    snl_aoi012x1 \ALUIS/U136  ( .ZN(\ALUIS/n3715 ), .A(\pgldi[12] ), .B(
        srcbsel), .C(allfbsel) );
    snl_oai222x0 \REGF/U471  ( .ZN(\REGF/RI_DPR[22] ), .A(\REGF/n8163 ), .B(
        \REGF/n8160 ), .C(\REGF/n8164 ), .D(\REGF/n8162 ), .E(\REGF/n8084 ), 
        .F(\REGF/n8151 ) );
    snl_invx05 \REGF/U741  ( .ZN(\REGF/n8145 ), .A(\pgldi[1] ) );
    snl_invx05 \REGF/U766  ( .ZN(\REGF/n8168 ), .A(\pgsdprlh[20] ) );
    snl_nand12x1 \ADOSEL/U61  ( .ZN(\ADOSEL/n4137 ), .A(\ADOSEL/n4157 ), .B(
        ph_word32_h) );
    snl_nand02x1 \ADOSEL/U46  ( .ZN(\ADOSEL/n4089 ), .A(ph_word32_h), .B(
        \ADOSEL/n4155 ) );
    snl_nand02x1 \PDOSEL/U150  ( .ZN(\PDOSEL/n124 ), .A(CDIN[20]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \REGF/U803  ( .ZN(\REGF/n8146 ), .A(\pkdptout[1] ) );
    snl_and02x1 \LDCHK/U97  ( .Z(\LDCHK/n3277 ), .A(\pgsadrh[1] ), .B(
        ph_word32_h) );
    snl_or04x1 \REGF/U818  ( .Z(\REGF/n8240 ), .A(\REGF/RO_ACC[19] ), .B(
        \REGF/RO_ACC[15] ), .C(\REGF/RO_ACC[28] ), .D(\REGF/RO_ACC[29] ) );
    snl_ao01b2x0 \RSTGN/U18  ( .Z(phrstihb), .A(\RSTGN/CRST_2H ), .B(
        \RSTGN/WRST_2H ), .C(phtri) );
    snl_and03x1 \RSTGN/U19  ( .Z(\RSTGN/n_6 ), .A(\RSTGN/WRST_1H ), .B(
        phrstith), .C(pgrstith) );
    snl_ffqx1 \RSTGN/CRST_1H_reg  ( .Q(\RSTGN/CRST_1H ), .D(CRST), .CP(SCLK)
         );
    snl_oai2222x0 \REGF/U360  ( .ZN(\REGF/RI_SRA12M[12] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8114 ), .C(\REGF/n8112 ), .D(\REGF/n8051 ), .E(\REGF/n8183 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8184 ) );
    snl_ao222x1 \CODEIF/U206  ( .Z(\CODEIF/n3853 ), .A(PA[15]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[12] ), .E(cif_byte), .F(PDLIN[12]
        ) );
    snl_muxi21x1 \CONS/U277  ( .ZN(\CONS/n538 ), .A(\CONS/n647 ), .B(
        \CONS/n641 ), .S(pk_pcser_h) );
    snl_oai122x0 \CODEIF/U221  ( .ZN(\CODEIF/pfctr415[0] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3865 ), .C(\CODEIF/n3866 ), .D(\CODEIF/n3867 ), .E(
        \CODEIF/n3868 ) );
    snl_xnor2x0 \CODEIF/U396  ( .ZN(\CODEIF/n3991 ), .A(CDIN[13]), .B(CDIN[14]
        ) );
    snl_xor2x0 \CODEIF/U417  ( .Z(\CODEIF/n4042 ), .A(\CODEIF/n4012 ), .B(
        \CODEIF/n4008 ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[0]  ( .Q(\pgld32[0] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[0] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_invx05 \LBUS/U630  ( .ZN(\LBUS/n1599 ), .A(pgadrovfh) );
    snl_nor02x1 \LBUS/U617  ( .ZN(\LBUS/n1592 ), .A(\LBUS/n1461 ), .B(
        \LBUS/n1593 ) );
    snl_nor04x0 \CONS/U147  ( .ZN(\CONS/n534 ), .A(\CONS/n710 ), .B(
        \CONS/n609 ), .C(\CONS/n607 ), .D(\CONS/n608 ) );
    snl_invx05 \PDOSEL/U94  ( .ZN(\PDOSEL/n77 ), .A(CDIN[33]) );
    snl_and08x1 \CONS/U160  ( .Z(\CONS/n345 ), .A(\CONS/n739 ), .B(\CONS/n740 
        ), .C(\CONS/n741 ), .D(\CONS/n742 ), .E(\CONS/n743 ), .F(\CONS/n744 ), 
        .G(\CONS/n745 ), .H(\CONS/n738 ) );
    snl_xnor2x0 \CONS/U250  ( .ZN(\CONS/n727 ), .A(\pk_idcx_h[17] ), .B(
        \pk_indx_h[17] ) );
    snl_nand02x1 \ALUIS/U44  ( .ZN(\pgaluina[28] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3686 ) );
    snl_xnor2x0 \LDCHK/U108  ( .ZN(\LDCHK/n3285 ), .A(\pgmuxout[16] ), .B(
        \pgmuxout[19] ) );
    snl_and02x1 \UPIF/U16  ( .Z(\ph_pdis_h[1] ), .A(\pk_rread_h[62] ), .B(
        \UPIF/n1046 ) );
    snl_nand02x2 \REGF/U385  ( .ZN(\REGF/n8230 ), .A(ph_oprtrs_h), .B(
        \REGF/n8228 ) );
    snl_invx2 \REGF/U404  ( .ZN(\REGF/n8217 ), .A(\ph_pdis_h[0] ) );
    snl_ao022x1 \REGF/U423  ( .Z(\REGF/RI_PCOH[10] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[10]), .C(\stream4[42] ), .D(\REGF/n8053 ) );
    snl_ao2222x1 \REGF/U538  ( .Z(\REGF/RI_SRDA[19] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[19]), .C(\pgldi[19] ), .D(\REGF/n8210 ), .E(\stream3[19] ), .F(
        \REGF/n8211 ), .G(\pkdptout[19] ), .H(\REGF/n8212 ) );
    snl_ao2222x1 \REGF/U556  ( .Z(\REGF/RI_SRDA[1] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[1]), .C(\pgldi[1] ), .D(\REGF/n8210 ), .E(\stream3[1] ), .F(
        \REGF/n8211 ), .G(\pkdptout[1] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U571  ( .ZN(\REGF/RI_ACC[30] ), .A(\REGF/n8060 ), .B(
        \REGF/n8215 ), .C(\REGF/n8061 ), .D(\REGF/n8216 ), .E(\REGF/n8062 ), 
        .F(\REGF/n8217 ) );
    snl_oai022x1 \REGF/U641  ( .ZN(\REGF/RI_TBAI[16] ), .A(\REGF/n8225 ), .B(
        \REGF/n8090 ), .C(\REGF/n8226 ), .D(\REGF/n8167 ) );
    snl_invx05 \REGF/U666  ( .ZN(\REGF/n8187 ), .A(\pgregadrh[10] ) );
    snl_oai012x1 \MAIN/U135  ( .A(ph_exstga_h), .B(\MAIN/n3618 ), .C(
        \MAIN/n3619 ) );
    snl_xor2x0 \CONS/U49  ( .Z(\CONS/n571 ), .A(\pk_saco_lh[20] ), .B(
        \pgsdprlh[20] ) );
    snl_oai012x1 \PDOSEL/U38  ( .ZN(PDH[54]), .A(\PDOSEL/n108 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nand02x1 \ADOSEL/U105  ( .ZN(\ADOSEL/n4139 ), .A(\pgbluext[16] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U63  ( .ZN(\pgaluinb[15] ), .A(\ALUIS/n3720 ), .B(
        \ALUIS/n3721 ) );
    snl_or03x1 \UPIF/U8  ( .Z(\UPIF/alusfterr ), .A(pkaluovf), .B(pkshterr), 
        .C(ph_lmterr_h) );
    snl_sffqenx1 \BLU/SRC_DATA_reg  ( .Q(pk_bitdatah), .D(1'b0), .EN(1'b1), 
        .SD(\BLU/SRC_DATA_M ), .SE(ph_bnolt_h), .CP(SCLK) );
    snl_oai222x0 \REGF/U608  ( .ZN(\REGF/RI_SPR[21] ), .A(\REGF/n8165 ), .B(
        \REGF/n8220 ), .C(\REGF/n8166 ), .D(\REGF/n8221 ), .E(\REGF/n8087 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U798  ( .ZN(\REGF/n8077 ), .A(\pkdptout[24] ) );
    snl_ao022x1 \BLUOS/U14  ( .Z(\pgbluext[26] ), .A(\pkbludgh[10] ), .B(
        ph_bit_h), .C(\pkdptout[10] ), .D(ph_word16_h) );
    snl_oai012x1 \LDIS/U132  ( .ZN(\pgldi[18] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3118 ), .C(\LDIS/n3115 ) );
    snl_or02x1 \CMPX/U23  ( .Z(\CMPX/n1051 ), .A(ph_sprsel2_h), .B(
        ph_dprsel2_h) );
    snl_xnor2x0 \CONS/U185  ( .ZN(\CONS/n665 ), .A(\pk_saco_lh[0] ), .B(
        \pgsdprlh[0] ) );
    snl_oai112x0 \PDOSEL/U56  ( .ZN(PDLOUT[12]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n98 ), .C(\PDOSEL/n136 ), .D(\PDOSEL/n137 ) );
    snl_mux21x1 \ALUSHT/U41  ( .Z(\pkdptout[11] ), .A(\ALUSHT/pkshtout[11] ), 
        .B(\ALUSHT/pkaluout[11] ), .S(\ALUSHT/n3112 ) );
    snl_nand02x1 \CODEIF/U354  ( .ZN(\CODEIF/n3904 ), .A(\CODEIF/pgctrinc[12] 
        ), .B(\CODEIF/n3945 ) );
    snl_invx05 \LDIS/U202  ( .ZN(\LDIS/n3146 ), .A(LIN[19]) );
    snl_nor04x0 \BLU/U323  ( .ZN(\BLU/n1487 ), .A(\BLU/n1530 ), .B(\BLU/n1528 
        ), .C(\BLU/n1531 ), .D(\BLU/n1532 ) );
    snl_nand02x1 \ALUIS/U164  ( .ZN(\ALUIS/n3659 ), .A(\pk_ada_h[1] ), .B(
        po_arsel_h) );
    snl_invx05 \REGF/U683  ( .ZN(\REGF/n8157 ), .A(PDLIN[28]) );
    snl_nor06x1 \REGF/U713  ( .ZN(\REGF/n8211 ), .A(ph_bdstenh), .B(ph_wdstenh
        ), .C(\REGF/n8233 ), .D(ph_wdsrdaselh), .E(\ph_pdis_h[9] ), .F(
        ph_btsrdaselh) );
    snl_xnor2x0 \CODEIF/U373  ( .ZN(\CODEIF/n3967 ), .A(CDIN[50]), .B(CDIN[47]
        ) );
    snl_invx05 \LDIS/U225  ( .ZN(\LDIS/n3151 ), .A(LIN[15]) );
    snl_aoi022x1 \ALUIS/U143  ( .ZN(\ALUIS/n3690 ), .A(\stream4[0] ), .B(
        immbsel), .C(\pk_adb_h[0] ), .D(po_brsel_h) );
    snl_xor2x0 \LDCHK/U69  ( .Z(\LDCHK/n3299 ), .A(\pgld32[12] ), .B(
        \pgld32[9] ) );
    snl_ao022x1 \LDIS/U115  ( .Z(\pgld16[8] ), .A(ph_selldl), .B(\pgld32[8] ), 
        .C(ph_selldh), .D(\pgld32[24] ) );
    snl_ao112x1 \PDOSEL/U71  ( .Z(PDLOUT[30]), .A(CDIN[30]), .B(\PDOSEL/n119 ), 
        .C(\pk_pdo_h[30] ), .D(\ph_cpudout[30] ) );
    snl_oai022x1 \BLU/U304  ( .ZN(\pkbludgh[12] ), .A(\BLU/n1464 ), .B(
        \BLU/n1474 ), .C(\BLU/n1475 ), .D(\BLU/n1476 ) );
    snl_invx05 \SAEXE/U142  ( .ZN(ph_trsc_h), .A(\SAEXE/n412 ) );
    snl_oai122x0 \ADOSEL/U14  ( .ZN(\pgmuxout[3] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4098 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4099 ), .E(
        \ADOSEL/n4100 ) );
    snl_invx05 \LBUS/U679  ( .ZN(\LBUS/n1444 ), .A(\LBUS/n1594 ) );
    snl_invx05 \PDOSEL/U102  ( .ZN(\PDOSEL/n98 ), .A(CDIN[44]) );
    snl_oai222x0 \REGF/U594  ( .ZN(\REGF/RI_ACC[7] ), .A(\REGF/n8127 ), .B(
        \REGF/n8215 ), .C(\REGF/n8128 ), .D(\REGF/n8216 ), .E(\REGF/n8129 ), 
        .F(\REGF/n8217 ) );
    snl_aoi012x1 \ALUIS/U86  ( .ZN(\ALUIS/n3703 ), .A(\pgldi[6] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_invx05 \BLU/U429  ( .ZN(\BLU/n1553 ), .A(\BLU/n1556 ) );
    snl_invx1 \REGF/U397  ( .ZN(\REGF/n8225 ), .A(\ph_pdis_h[10] ) );
    snl_ao022x1 \REGF/U416  ( .Z(\REGF/RI_PCOH[17] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[17]), .C(\stream4[49] ), .D(\REGF/n8053 ) );
    snl_ao022x1 \REGF/U431  ( .Z(\REGF/RI_PCOH[2] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[2]), .C(\stream4[34] ), .D(\REGF/n8053 ) );
    snl_invx05 \REGF/U691  ( .ZN(\REGF/n8087 ), .A(PDLIN[21]) );
    snl_invx05 \REGF/U734  ( .ZN(\REGF/n8075 ), .A(PDLIN[25]) );
    snl_invx05 \CODEIF/U268  ( .ZN(\CODEIF/n3872 ), .A(\CODEIF/pfctr[2] ) );
    snl_xnor2x0 \CONS/U219  ( .ZN(\CONS/n704 ), .A(\pk_idcz_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[14]  ( .Q(\ph_segset_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[14]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_and02x1 \REG_2/U148  ( .Z(\ph_cpudout[18] ), .A(\ph_segset_h[18] ), 
        .B(seg_cnfg_h) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[27]  ( .Q(\ph_segset_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[27]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_oai122x0 \ADOSEL/U33  ( .ZN(\pgmuxout[22] ), .A(\ADOSEL/n4108 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4107 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4145 ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[10]  ( .Q(\pgld32[10] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexcl[10] ), .SE(lo_data_lth), .CP(SCLK
        ) );
    snl_ao022x1 \CMPX/U6  ( .Z(ph_bitsrc_h), .A(ph_bitsrch), .B(ph_saexe_sth), 
        .C(po_bitsrc_h), .D(\CMPX/n1047 ) );
    snl_nor02x1 \PDOSEL/U125  ( .ZN(\PDOSEL/n161 ), .A(\ph_cpudout[18] ), .B(
        \pk_pdo_h[18] ) );
    snl_nor02x1 \CONS/U129  ( .ZN(\CONS/n667 ), .A(\CONS/n576 ), .B(
        \CONS/n577 ) );
    snl_xor2x0 \CONS/U99  ( .Z(\CONS/n617 ), .A(\pk_idcy_h[18] ), .B(
        \pk_indy_h[18] ) );
    snl_invx05 \REGF/U701  ( .ZN(\REGF/n8102 ), .A(PDLIN[16]) );
    snl_nor02x1 \PDOSEL/U110  ( .ZN(\PDOSEL/n157 ), .A(\ph_cpudout[6] ), .B(
        \pk_pdo_h[6] ) );
    snl_aoi012x1 \ALUIS/U94  ( .ZN(\ALUIS/n3753 ), .A(\pgldi[31] ), .B(srcbsel
        ), .C(allfbsel) );
    snl_oai222x0 \REGF/U586  ( .ZN(\REGF/RI_ACC[15] ), .A(\REGF/n8103 ), .B(
        \REGF/n8215 ), .C(\REGF/n8104 ), .D(\REGF/n8216 ), .E(\REGF/n8105 ), 
        .F(\REGF/n8217 ) );
    snl_ffqsnx1 \LBUS/l_wr_reg  ( .Q(LWR), .D(phrstith), .SN(n10734), .CP(SCLK
        ) );
    snl_ffandx1 \RSTGN/WRST_2H_reg  ( .Q(\RSTGN/WRST_2H ), .A(CRWE), .B(
        \RSTGN/n_6 ), .CP(SCLK) );
    snl_oai2222x0 \REGF/U355  ( .ZN(\REGF/RI_SRA12M[20] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8090 ), .C(\REGF/n8088 ), .D(\REGF/n8051 ), .E(\REGF/n8167 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8168 ) );
    snl_oai022x1 \REGF/U372  ( .ZN(\REGF/RI_TBAI[11] ), .A(\REGF/n8225 ), .B(
        \REGF/n8105 ), .C(\REGF/n8226 ), .D(\REGF/n8177 ) );
    snl_and02x1 \REGF/U563  ( .Z(\REGF/RO_LPSAS2156[5] ), .A(ph_sastlth), .B(
        \REGF/RO_EST1[7] ) );
    snl_invx05 \REGF/U726  ( .ZN(\REGF/n8144 ), .A(PDLIN[2]) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[6]  ( .Q(\REGF/RO_LLPSAS[8] ), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[6] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_oai122x0 \ADOSEL/U21  ( .ZN(\pgmuxout[10] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4119 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4120 ), .E(
        \ADOSEL/n4121 ) );
    snl_nand02x1 \PDOSEL/U137  ( .ZN(\PDOSEL/n146 ), .A(CDIN[7]), .B(
        \PDOSEL/n119 ) );
    snl_nand02x1 \CODEIF/U346  ( .ZN(\CODEIF/n3874 ), .A(\CODEIF/pgctrinc[2] ), 
        .B(\CODEIF/n3945 ) );
    snl_invx05 \MAIN/U149  ( .ZN(\MAIN/n3628 ), .A(\MAIN/ph_rdwr2selh ) );
    snl_ao022x1 \LDIS/U120  ( .Z(\pgldi[11] ), .A(ph_word32_h), .B(
        \pgld32[11] ), .C(\pgld16[11] ), .D(ph_word16_h) );
    snl_sffqensnx2 \REG_2/ph_retcnt_h_reg[1]  ( .Q(\REG_2/ph_retcnt_h[1] ), 
        .D(1'b0), .EN(1'b1), .SN(\REG_2/n435 ), .SD(PDLIN[1]), .SE(ret_cont_wr
        ), .CP(SCLK) );
    snl_xnor2x0 \CONS/U197  ( .ZN(\CONS/n677 ), .A(\pk_pc_h[14] ), .B(
        \pk_pcs2_h[14] ) );
    snl_oai112x0 \PDOSEL/U44  ( .ZN(PDLOUT[10]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n96 ), .C(\PDOSEL/n115 ), .D(\PDOSEL/n116 ) );
    snl_invx05 \LDIS/U210  ( .ZN(\LDIS/n3138 ), .A(LIN[23]) );
    snl_nor02x1 \BLU/U331  ( .ZN(\BLU/n1466 ), .A(\BLU/n1544 ), .B(\BLU/n1545 
        ) );
    snl_xor2x0 \CODEIF/U361  ( .Z(\CODEIF/n4022 ), .A(\CODEIF/n4023 ), .B(
        \CODEIF/n3999 ) );
    snl_oai022x1 \BLU/U316  ( .ZN(\pkbludgh[0] ), .A(\BLU/n1464 ), .B(
        \BLU/n1510 ), .C(\BLU/n1511 ), .D(\BLU/n1512 ) );
    snl_nand02x1 \ALUIS/U38  ( .ZN(\pgaluina[22] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3680 ) );
    snl_nand02x1 \ALUIS/U56  ( .ZN(\pgaluinb[8] ), .A(\ALUIS/n3706 ), .B(
        \ALUIS/n3707 ) );
    snl_nand02x1 \ALUIS/U151  ( .ZN(\ALUIS/n3689 ), .A(\pk_ada_h[31] ), .B(
        po_arsel_h) );
    snl_ao022x1 \BLUOS/U21  ( .Z(\pgbluext[2] ), .A(\pkbludgh[2] ), .B(
        ph_bit_h), .C(\pkdptout[2] ), .D(ph_word16_h) );
    snl_ao022x1 \LDIS/U107  ( .Z(\pgld16[4] ), .A(ph_selldl), .B(\pgld32[4] ), 
        .C(ph_selldh), .D(\pgld32[20] ) );
    snl_nor02x1 \CMPX/U16  ( .ZN(ph_adrdec_h), .A(\CMPX/n1047 ), .B(
        \CMPX/n1050 ) );
    snl_ffqrnx1 \LBUS/ilt_reg[5]  ( .Q(\LBUS/ilt[5] ), .D(\LBUS/nlt[5] ), .RN(
        n10734), .CP(SCLK) );
    snl_aoi012x1 \CONS/U35  ( .ZN(\CONS/n543 ), .A(word32odtrh), .B(
        \CONS/n544 ), .C(\CONS/n540 ) );
    snl_oai112x0 \PDOSEL/U63  ( .ZN(PDLOUT[16]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n102 ), .C(\PDOSEL/n150 ), .D(\PDOSEL/n151 ) );
    snl_nand13x1 \BLU/U378  ( .ZN(\BLU/n1540 ), .A(\BLU/n1533 ), .B(
        \BLU/n1489 ), .C(\BLU/n1572 ) );
    snl_ffqrnx1 \SAEXE/ph_lber1_h_reg  ( .Q(\SAEXE/ph_lber1_h ), .D(ph_lberr), 
        .RN(n10735), .CP(SCLK) );
    snl_oai022x1 \REGF/U653  ( .ZN(\REGF/RI_TBAI[1] ), .A(\REGF/n8225 ), .B(
        \REGF/n8135 ), .C(\REGF/n8226 ), .D(\REGF/n8197 ) );
    snl_muxi21x1 \LDIS/U169  ( .ZN(\LDIS/ldexcl[3] ), .A(\LDIS/n3145 ), .B(
        \LDIS/n3146 ), .S(\LDIS/n3134 ) );
    snl_oa112x1 \LBUS/U599  ( .Z(\LBUS/n1448 ), .A(\LBUS/n1452 ), .B(
        \LBUS/ilt[2] ), .C(\LBUS/n1453 ), .D(\LBUS/n1430 ) );
    snl_invx05 \REGF/U674  ( .ZN(\REGF/n8195 ), .A(\pgregadrh[6] ) );
    snl_ao013x1 \MAIN/U127  ( .Z(ph_stage_ah), .A(\MAIN/n3618 ), .B(
        \MAIN/n3619 ), .C(stage_a), .D(ph_exstga_h) );
    snl_nor02x1 \LDCHK/U32  ( .ZN(LPOUT[1]), .A(\LDCHK/n3231 ), .B(
        \LDCHK/n3233 ) );
    snl_nor02x1 \SAEXE/U119  ( .ZN(\SAEXE/n416 ), .A(ph_lblockh), .B(
        \SAEXE/n423 ) );
    snl_xor2x0 \CODEIF/U328  ( .Z(\CODEIF/n4007 ), .A(CDOUT[33]), .B(CDOUT[31]
        ) );
    snl_nand02x1 \ALUIS/U71  ( .ZN(\pgaluinb[23] ), .A(\ALUIS/n3736 ), .B(
        \ALUIS/n3737 ) );
    snl_aoi012x1 \ALUIS/U118  ( .ZN(\ALUIS/n3731 ), .A(\pgldi[20] ), .B(
        srcbsel), .C(allfbsel) );
    snl_oai222x0 \REGF/U444  ( .ZN(\REGF/RI_EACC[21] ), .A(\REGF/n8085 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8086 ), .E(\REGF/n8087 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U478  ( .ZN(\REGF/RI_DPR[15] ), .A(\REGF/n8177 ), .B(
        \REGF/n8160 ), .C(\REGF/n8178 ), .D(\REGF/n8162 ), .E(\REGF/n8105 ), 
        .F(\REGF/n8151 ) );
    snl_ao2222x1 \REGF/U544  ( .Z(\REGF/RI_SRDA[13] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[13]), .C(\pgldi[13] ), .D(\REGF/n8210 ), .E(\stream3[13] ), .F(
        \REGF/n8211 ), .G(\pkdptout[13] ), .H(\REGF/n8212 ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[23]  ( .Q(\pgld32[23] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[23] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[19]  ( .Q(\ph_segset_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[19]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_invx05 \REGF/U748  ( .ZN(\REGF/n8109 ), .A(\pgldi[13] ) );
    snl_invx1 \CODEIF/U214  ( .ZN(\CODEIF/n3861 ), .A(\CODEIF/n3860 ) );
    snl_xor2x0 \CODEIF/U384  ( .Z(\CODEIF/n3934 ), .A(\CODEIF/n3979 ), .B(
        \CODEIF/n4032 ) );
    snl_ao022x1 \REG_2/U134  ( .Z(\ph_cpudout[4] ), .A(\ph_segset_h[4] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[4] ), .D(ret_cont_h) );
    snl_xor2x0 \CODEIF/U405  ( .Z(\CODEIF/n4038 ), .A(\CODEIF/n3998 ), .B(
        \CODEIF/n3994 ) );
    snl_xnor2x0 \CONS/U265  ( .ZN(\CONS/n739 ), .A(\pk_idcw_h[21] ), .B(
        \pk_indw_h[21] ) );
    snl_invx05 \ADOSEL/U68  ( .ZN(\ADOSEL/n4096 ), .A(\pkdptout[2] ) );
    snl_nor03x0 \LBUS/U605  ( .ZN(ph_lpdilth), .A(LDS), .B(ph_lbwrh), .C(
        \LBUS/n1425 ) );
    snl_invx05 \LBUS/U622  ( .ZN(\LBUS/n1417 ), .A(ph_tirtendh) );
    snl_sffqenrnx1 \LBUS/ph_exstga_h_reg  ( .Q(ph_exstga_h), .D(1'b0), .EN(
        1'b1), .RN(n10734), .SD(\LBUS/*cell*3982/U70/CONTROL1 ), .SE(
        \LBUS/*cell*3982/U200/CONTROL1 ), .CP(SCLK) );
    snl_and08x1 \CONS/U155  ( .Z(\CONS/n519 ), .A(\CONS/n727 ), .B(\CONS/n728 
        ), .C(\CONS/n729 ), .D(\CONS/n730 ), .E(\CONS/n731 ), .F(\CONS/n732 ), 
        .G(\CONS/n733 ), .H(\CONS/n726 ) );
    snl_invx05 \PDOSEL/U86  ( .ZN(\PDOSEL/n113 ), .A(CDIN[59]) );
    snl_nand02x1 \PDOSEL/U159  ( .ZN(\PDOSEL/n122 ), .A(CDIN[13]), .B(
        \PDOSEL/n119 ) );
    snl_oai122x0 \CODEIF/U228  ( .ZN(\CODEIF/pfctr415[7] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3887 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3888 ), .E(
        \CODEIF/n3889 ) );
    snl_oai122x0 \CODEIF/U233  ( .ZN(\CODEIF/pfctr415[12] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3902 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3903 ), .E(
        \CODEIF/n3904 ) );
    snl_sffqenrnx1 \MAIN/ph_lmterrh_reg  ( .Q(phlmterrh), .D(1'b0), .EN(1'b1), 
        .RN(\MAIN/n3611 ), .SD(\MAIN/*cell*4603/U1/CONTROL1 ), .SE(
        \MAIN/*cell*4603/U15/CONTROL1 ), .CP(SCLK) );
    snl_xnor2x0 \CONS/U172  ( .ZN(\CONS/n649 ), .A(\pgsdprlh[14] ), .B(
        \pk_saco_lh[14] ) );
    snl_xor2x0 \CODEIF/U422  ( .Z(\CODEIF/n4029 ), .A(\CODEIF/n4043 ), .B(
        CDOUT[10]) );
    snl_xnor2x0 \CONS/U242  ( .ZN(\CONS/n525 ), .A(\pk_idcy_h[7] ), .B(
        \pk_indy_h[7] ) );
    snl_xnor2x0 \CONS/U259  ( .ZN(\CONS/n346 ), .A(\pk_idcx_h[6] ), .B(
        \pk_indx_h[6] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[10]  ( .Q(\ph_segset_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[10]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_invx05 \REGF/U753  ( .ZN(\REGF/n8190 ), .A(\pgsdprlh[9] ) );
    snl_invx05 \REGF/U774  ( .ZN(\REGF/n8180 ), .A(\pgsdprlh[14] ) );
    snl_sffqenrnx1 \REGF/RO_LPSAS_reg[11]  ( .Q(\REGF/RO_LLPSAS[15] ), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/n8052 ), .SD(\REGF/RO_LPSAS2156[11] ), .SE(
        \REGF/n_2734 ), .CP(SCLK) );
    snl_xnor2x0 \CONS/U169  ( .ZN(\CONS/n555 ), .A(\pk_saco_hh[31] ), .B(
        \pgsdprhh[31] ) );
    snl_invx05 \ADOSEL/U73  ( .ZN(\ADOSEL/n4123 ), .A(\pkdptout[11] ) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[14]  ( .Q(\pgld32[14] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexcl[14] ), .SE(lo_data_lth), .CP(SCLK
        ) );
    snl_invx05 \ADOSEL/U54  ( .ZN(\ADOSEL/n4104 ), .A(\pkdptout[21] ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[23]  ( .Q(\ph_segset_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[23]), .SE(seg_config_wr
        ), .CP(SCLK) );
    snl_or04x1 \LDCHK/U85  ( .Z(\LDCHK/n3309 ), .A(\pgld32[9] ), .B(
        \pgld32[28] ), .C(\pgld32[21] ), .D(\pgld32[12] ) );
    snl_oai113x0 \LBUS/U639  ( .ZN(\LBUS/n1434 ), .A(\LBUS/n1602 ), .B(
        \LBUS/n1597 ), .C(\LBUS/n1406 ), .D(\LBUS/n1432 ), .E(\LBUS/n1428 ) );
    snl_nand02x1 \PDOSEL/U142  ( .ZN(\PDOSEL/n144 ), .A(CDIN[2]), .B(
        \PDOSEL/n119 ) );
    snl_oai2222x0 \REGF/U369  ( .ZN(\REGF/RI_SRA12M[0] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8150 ), .C(\REGF/n8148 ), .D(\REGF/n8051 ), .E(\REGF/n8229 ), 
        .F(\REGF/n8207 ), .G(\REGF/n8230 ), .H(\REGF/n8208 ) );
    snl_oai222x0 \REGF/U463  ( .ZN(\REGF/RI_EACC[2] ), .A(\REGF/n8142 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8143 ), .E(\REGF/n8144 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U578  ( .ZN(\REGF/RI_ACC[23] ), .A(\REGF/n8079 ), .B(
        \REGF/n8215 ), .C(\REGF/n8080 ), .D(\REGF/n8216 ), .E(\REGF/n8081 ), 
        .F(\REGF/n8217 ) );
    snl_oai022x1 \REGF/U648  ( .ZN(\REGF/RI_TBAI[6] ), .A(\REGF/n8225 ), .B(
        \REGF/n8120 ), .C(\REGF/n8226 ), .D(\REGF/n8187 ) );
    snl_invx05 \REGF/U811  ( .ZN(\REGF/n8113 ), .A(\pkdptout[12] ) );
    snl_xor2x0 \CODEIF/U333  ( .Z(\CODEIF/n4014 ), .A(CDOUT[15]), .B(CDOUT[16]
        ) );
    snl_invx05 \BLU/U344  ( .ZN(\BLU/n1559 ), .A(\pgbitnoh[3] ) );
    snl_aoi022x1 \ALUIS/U103  ( .ZN(\ALUIS/n3746 ), .A(\stream4[28] ), .B(
        immbsel), .C(\pk_adb_h[28] ), .D(po_brsel_h) );
    snl_invx05 \LDIS/U155  ( .ZN(\LDIS/n3130 ), .A(\pgld32[30] ) );
    snl_mux21x1 \ALUSHT/U26  ( .Z(\pkdptout[25] ), .A(\ALUSHT/pkshtout[25] ), 
        .B(\ALUSHT/pkaluout[25] ), .S(\ALUSHT/n3112 ) );
    snl_aoi022x1 \CONS/U67  ( .ZN(\CONS/n584 ), .A(\CONS/n551 ), .B(
        \CONS/n585 ), .C(\pgsdprlh[4] ), .D(\CONS/SACO[0] ) );
    snl_nand12x1 \SAEXE/U102  ( .ZN(\SAEXE/*cell*3651/U11/CONTROL1 ), .A(
        \pk_rwrit_h[49] ), .B(\SAEXE/n412 ) );
    snl_aoi022x1 \LBUS/U695  ( .ZN(\LBUS/n1418 ), .A(ph_byrtendh), .B(
        \LBUS/ph_lbusylth ), .C(\LBUS/n1604 ), .D(\LBUS/n1459 ) );
    snl_oai012x1 \PDOSEL/U31  ( .ZN(PDH[47]), .A(\PDOSEL/n101 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_invx05 \SAEXE/U125  ( .ZN(\SAEXE/n413 ), .A(ph_saexe_sth) );
    snl_xnor2x0 \LDCHK/U101  ( .ZN(\LDCHK/n3278 ), .A(\pgmuxout[26] ), .B(
        \pgmuxout[29] ) );
    snl_muxi21x1 \LDIS/U172  ( .ZN(\LDIS/ldexcl[15] ), .A(\LDIS/n3151 ), .B(
        \LDIS/n3152 ), .S(\LDIS/n3134 ) );
    snl_sffqenrnx1 \LDIS/pgld32h_reg[19]  ( .Q(\pgld32[19] ), .D(1'b0), .EN(
        1'b1), .RN(n10736), .SD(\LDIS/ldexch[19] ), .SE(up_data_lth), .CP(SCLK
        ) );
    snl_nand04x0 \CONS/U40  ( .ZN(\CONS/n552 ), .A(\CONS/n553 ), .B(
        \CONS/n554 ), .C(\CONS/n555 ), .D(\CONS/n556 ) );
    snl_oai012x1 \PDOSEL/U16  ( .ZN(PDH[32]), .A(\PDOSEL/n74 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_oai012x1 \LBUS/U582  ( .ZN(ph_d76lth), .A(\LBUS/n1444 ), .B(
        \LBUS/n1445 ), .C(\LBUS/n1446 ) );
    snl_oai222x0 \REGF/U486  ( .ZN(\REGF/RI_DPR[7] ), .A(\REGF/n8193 ), .B(
        \REGF/n8160 ), .C(\REGF/n8194 ), .D(\REGF/n8162 ), .E(\REGF/n8129 ), 
        .F(\REGF/n8151 ) );
    snl_oai222x0 \REGF/U626  ( .ZN(\REGF/RI_SPR[3] ), .A(\REGF/n8201 ), .B(
        \REGF/n8220 ), .C(\REGF/n8202 ), .D(\REGF/n8221 ), .E(\REGF/n8141 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \CODEIF/U284  ( .ZN(\CODEIF/n3902 ), .A(\CODEIF/pfctr[12] ) );
    snl_xor2x0 \CODEIF/U314  ( .Z(\CODEIF/n3958 ), .A(\CODEIF/n3987 ), .B(
        \CODEIF/n3988 ) );
    snl_aoi012x1 \ALUIS/U124  ( .ZN(\ALUIS/n3727 ), .A(\pgldi[18] ), .B(
        srcbsel), .C(allfbsel) );
    snl_xor2x0 \LDCHK/U60  ( .Z(\LDCHK/n3260 ), .A(\LDCHK/n3286 ), .B(
        \LDCHK/n3287 ) );
    snl_nand02x1 \BLU/U363  ( .ZN(\BLU/n1483 ), .A(\BLU/n1570 ), .B(
        \BLU/n1562 ) );
    snl_invx05 \PDOSEL/U78  ( .ZN(\PDOSEL/n95 ), .A(CDIN[41]) );
    snl_ao022x1 \REGF/U516  ( .Z(\REGF/RI_PCOL[9] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[9]), .C(\REGF/n8209 ), .D(\stream4[9] ) );
    snl_ao2222x1 \REGF/U531  ( .Z(\REGF/RI_SRDA[26] ), .A(PDLIN[26]), .B(
        \ph_pdis_h[9] ), .C(\pgldi[26] ), .D(\REGF/n8210 ), .E(\stream3[26] ), 
        .F(\REGF/n8211 ), .G(\pkdptout[26] ), .H(\REGF/n8212 ) );
    snl_nand02x2 \ALUIS/U23  ( .ZN(\pgaluina[9] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3667 ) );
    snl_oai222x0 \REGF/U601  ( .ZN(\REGF/RI_ACC[0] ), .A(\REGF/n8148 ), .B(
        \REGF/n8215 ), .C(\REGF/n8149 ), .D(\REGF/n8216 ), .E(\REGF/n8150 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U791  ( .ZN(\REGF/n8061 ), .A(\pkdptout[30] ) );
    snl_nand02x1 \ADOSEL/U96  ( .ZN(\ADOSEL/n4147 ), .A(\pgbluext[8] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \MAIN/U152  ( .ZN(\MAIN/n3626 ), .A(pgadrovfh), .B(
        \MAIN/n3633 ) );
    snl_xor2x0 \LDCHK/U47  ( .Z(\LDCHK/n3232 ), .A(\LDCHK/n3262 ), .B(
        \LDCHK/n3263 ) );
    snl_invx05 \CODEIF/U261  ( .ZN(\CODEIF/n3885 ), .A(PDLIN[6]) );
    snl_invx05 \LDIS/U197  ( .ZN(\LDIS/n3149 ), .A(LIN[1]) );
    snl_nand02x1 \LBUS/U657  ( .ZN(\LBUS/n1413 ), .A(ph_ioselh), .B(ph_lbussth
        ) );
    snl_nand12x1 \CONS/U120  ( .ZN(\CONS/n639 ), .A(\pk_saseo_h[0] ), .B(
        \CONS/n640 ) );
    snl_xnor2x0 \CONS/U210  ( .ZN(\CONS/n692 ), .A(\pk_pc_h[18] ), .B(
        \pk_pcs1_h[18] ) );
    snl_oai013x0 \BLU/U407  ( .ZN(\BLU/n1578 ), .A(\BLU/n1555 ), .B(
        \poalufnc[1] ), .C(\poalufnc[0] ), .D(\BLU/n1579 ) );
    snl_and02x1 \REG_2/U141  ( .Z(\ph_cpudout[11] ), .A(\ph_segset_h[11] ), 
        .B(seg_cnfg_h) );
    snl_nand13x1 \BLU/U386  ( .ZN(\BLU/n1545 ), .A(\BLU/n1550 ), .B(
        \BLU/n1571 ), .C(\BLU/n1477 ) );
    snl_xor2x0 \CODEIF/U246  ( .Z(CPOUT[2]), .A(\CODEIF/n3938 ), .B(
        \CODEIF/n3939 ) );
    snl_nor02x1 \LBUS/U567  ( .ZN(ph_pdlen_h), .A(\LBUS/n1412 ), .B(
        \LBUS/n1391 ) );
    snl_xnor2x0 \CONS/U237  ( .ZN(\CONS/n724 ), .A(\pk_idcy_h[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \BLU/U420  ( .ZN(\BLU/n1535 ), .A(\BLU/n1495 ) );
    snl_oai2222x0 \REGF/U354  ( .ZN(\REGF/RI_SRA12M[21] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8087 ), .C(\REGF/n8085 ), .D(\REGF/n8051 ), .E(\REGF/n8165 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8166 ) );
    snl_oai2222x0 \REGF/U361  ( .ZN(\REGF/RI_SRA12M[10] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8120 ), .C(\REGF/n8118 ), .D(\REGF/n8051 ), .E(\REGF/n8187 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8188 ) );
    snl_oai2222x0 \REGF/U384  ( .ZN(\REGF/RI_SRA12M[7] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8129 ), .C(\REGF/n8127 ), .D(\REGF/n8051 ), .E(\REGF/n8193 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8194 ) );
    snl_ao022x1 \REGF/U422  ( .Z(\REGF/RI_PCOH[11] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[11]), .C(\stream4[43] ), .D(\REGF/n8053 ) );
    snl_ao2222x1 \REGF/U539  ( .Z(\REGF/RI_SRDA[18] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[18]), .C(\pgldi[18] ), .D(\REGF/n8210 ), .E(\stream3[18] ), .F(
        \REGF/n8211 ), .G(\pkdptout[18] ), .H(\REGF/n8212 ) );
    snl_oai222x0 \REGF/U609  ( .ZN(\REGF/RI_SPR[20] ), .A(\REGF/n8167 ), .B(
        \REGF/n8220 ), .C(\REGF/n8168 ), .D(\REGF/n8221 ), .E(\REGF/n8090 ), 
        .F(\REGF/n8218 ) );
    snl_ao022x1 \BLUOS/U15  ( .Z(\pgbluext[27] ), .A(\pkbludgh[11] ), .B(
        ph_bit_h), .C(\pkdptout[11] ), .D(ph_word16_h) );
    snl_sffqenrnx1 \LDIS/pgld32l_reg[4]  ( .Q(\pgld32[4] ), .D(1'b0), .EN(1'b1
        ), .RN(n10736), .SD(\LDIS/ldexcl[4] ), .SE(lo_data_lth), .CP(SCLK) );
    snl_ffqrnx1 \LBUS/access_en_h_reg  ( .Q(\LBUS/access_en_h ), .D(LASIN), 
        .RN(n10734), .CP(SCLK) );
    snl_xor2x0 \CONS/U107  ( .Z(\CONS/n625 ), .A(\pk_idcx_h[12] ), .B(
        \pk_indx_h[12] ) );
    snl_mux21x1 \ALUSHT/U40  ( .Z(\pkdptout[12] ), .A(\ALUSHT/pkshtout[12] ), 
        .B(\ALUSHT/pkaluout[12] ), .S(\ALUSHT/n3112 ) );
    snl_nor03x0 \LBUS/U670  ( .ZN(ph_d53lth), .A(LDS), .B(ph_byrtendh), .C(
        \LBUS/n1459 ) );
    snl_xor2x0 \CONS/U82  ( .Z(\CONS/n600 ), .A(\pk_pcs1_h[0] ), .B(
        \pk_pc_h[0] ) );
    snl_invx05 \REGF/U799  ( .ZN(\REGF/n8080 ), .A(\pkdptout[23] ) );
    snl_oai012x1 \LDIS/U133  ( .ZN(\pgldi[19] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3119 ), .C(\LDIS/n3115 ) );
    snl_ao022x1 \CMPX/U22  ( .Z(ph_sprtrs_h), .A(ph_sprsel2_h), .B(
        ph_saexe_sth), .C(po_sprtrs_h), .D(\CMPX/n1047 ) );
    snl_xnor2x0 \CONS/U184  ( .ZN(\CONS/n660 ), .A(\pgsdprlh[11] ), .B(
        \pk_saco_lh[11] ) );
    snl_oai112x0 \PDOSEL/U57  ( .ZN(PDLOUT[9]), .A(\PDOSEL/n95 ), .B(
        \PDOSEL/n114 ), .C(\PDOSEL/n138 ), .D(\PDOSEL/n139 ) );
    snl_invx05 \REGF/U682  ( .ZN(\REGF/n8158 ), .A(\pgsdprhh[28] ) );
    snl_ffqx1 \REGF/D2_DTFL_reg  ( .Q(\REGF/D2_DTFL ), .D(DTFL), .CP(SCLK) );
    snl_nand02x1 \CODEIF/U355  ( .ZN(\CODEIF/n3901 ), .A(\CODEIF/pgctrinc[11] 
        ), .B(\CODEIF/n3945 ) );
    snl_nand02x1 \ALUIS/U165  ( .ZN(\ALUIS/n3677 ), .A(\pk_ada_h[19] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U203  ( .ZN(\LDIS/n3143 ), .A(LIN[4]) );
    snl_nor02x1 \BLU/U322  ( .ZN(\BLU/n1484 ), .A(\BLU/n1528 ), .B(\BLU/n1529 
        ) );
    snl_oai122x0 \ADOSEL/U15  ( .ZN(\pgmuxout[4] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4101 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4102 ), .E(
        \ADOSEL/n4103 ) );
    snl_xnor2x0 \CODEIF/U372  ( .ZN(\CODEIF/n3965 ), .A(CDIN[56]), .B(CDIN[55]
        ) );
    snl_aoi012x1 \ALUIS/U142  ( .ZN(\ALUIS/n3691 ), .A(\pgldi[0] ), .B(srcbsel
        ), .C(allfbsel) );
    snl_invx05 \LDIS/U224  ( .ZN(\LDIS/n3154 ), .A(LIN[30]) );
    snl_oai022x1 \BLU/U305  ( .ZN(\pkbludgh[11] ), .A(\BLU/n1464 ), .B(
        \BLU/n1477 ), .C(\BLU/n1478 ), .D(\BLU/n1479 ) );
    snl_xor2x0 \LDCHK/U68  ( .Z(\LDCHK/n3298 ), .A(\pgld32[10] ), .B(
        \pgld32[13] ) );
    snl_oai022x1 \SAEXE/U143  ( .ZN(\SAEXE/n430 ), .A(\SAEXE/n423 ), .B(
        \SAEXE/n431 ), .C(\SAEXE/n427 ), .D(\SAEXE/n428 ) );
    snl_ao022x1 \LDIS/U114  ( .Z(\pgldi[8] ), .A(ph_word32_h), .B(\pgld32[8] ), 
        .C(\pgld16[8] ), .D(ph_word16_h) );
    snl_oai112x0 \PDOSEL/U70  ( .ZN(PDLOUT[5]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n81 ), .C(\PDOSEL/n162 ), .D(\PDOSEL/n163 ) );
    snl_invx05 \PDOSEL/U103  ( .ZN(\PDOSEL/n97 ), .A(CDIN[43]) );
    snl_and12x1 \REGF/U712  ( .Z(\REGF/n8212 ), .A(\ph_pdis_h[9] ), .B(
        ph_wdstenh) );
    snl_aoi022x1 \ALUIS/U87  ( .ZN(\ALUIS/n3702 ), .A(\stream4[6] ), .B(
        immbsel), .C(\pk_adb_h[6] ), .D(po_brsel_h) );
    snl_invx05 \LBUS/U678  ( .ZN(\LBUS/n1443 ), .A(\LBUS/n1592 ) );
    snl_invx05 \BLU/U428  ( .ZN(\BLU/n1549 ), .A(\BLU/n1465 ) );
    snl_invx05 \CODEIF/U269  ( .ZN(\CODEIF/n3873 ), .A(PDLIN[2]) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[5]  ( .Q(CA[5]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3846 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_xnor2x0 \CONS/U218  ( .ZN(\CONS/n708 ), .A(\pk_idcz_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_and02x1 \REG_2/U149  ( .Z(\ph_cpudout[19] ), .A(\ph_segset_h[19] ), 
        .B(seg_cnfg_h) );
    snl_or02x1 \REGF/U405  ( .Z(\REGF/n_2734 ), .A(\pk_rwrit_h[48] ), .B(
        ph_sastlth) );
    snl_oai222x0 \REGF/U570  ( .ZN(\REGF/RI_ACC[31] ), .A(\REGF/n8054 ), .B(
        \REGF/n8215 ), .C(\REGF/n8057 ), .D(\REGF/n8216 ), .E(\REGF/n8058 ), 
        .F(\REGF/n8217 ) );
    snl_oai222x0 \REGF/U595  ( .ZN(\REGF/RI_ACC[6] ), .A(\REGF/n8130 ), .B(
        \REGF/n8215 ), .C(\REGF/n8131 ), .D(\REGF/n8216 ), .E(\REGF/n8132 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U735  ( .ZN(\REGF/n8076 ), .A(\pgldi[24] ) );
    snl_oai122x0 \ADOSEL/U32  ( .ZN(\pgmuxout[21] ), .A(\ADOSEL/n4105 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4104 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4144 ) );
    snl_ao022x4 \CMPX/U7  ( .Z(ph_word16_h), .A(ph_word16h), .B(ph_saexe_sth), 
        .C(srctype1), .D(\CMPX/n1047 ) );
    snl_nor02x1 \PDOSEL/U124  ( .ZN(\PDOSEL/n131 ), .A(\pk_pdo_h[19] ), .B(
        \ph_cpudout[19] ) );
    snl_oai013x0 \CONS/U128  ( .ZN(\CONS/n638 ), .A(\CONS/n664 ), .B(
        \CONS/n574 ), .C(\CONS/n575 ), .D(\CONS/n540 ) );
    snl_or04x1 \REGF/U819  ( .Z(\REGF/n8241 ), .A(\REGF/RO_ACC[18] ), .B(
        \REGF/RO_ACC[21] ), .C(\REGF/RO_ACC[24] ), .D(\REGF/RO_ACC[16] ) );
    snl_ao222x1 \CODEIF/U207  ( .Z(\CODEIF/n3854 ), .A(PA[16]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[13] ), .E(cif_byte), .F(PDLIN[13]
        ) );
    snl_xnor2x0 \CODEIF/U397  ( .ZN(\CODEIF/n4035 ), .A(CDIN[4]), .B(CDIN[2])
         );
    snl_xor2x0 \CODEIF/U416  ( .Z(\CODEIF/n4027 ), .A(\CODEIF/n4041 ), .B(
        CDOUT[24]) );
    snl_muxi21x1 \CONS/U276  ( .ZN(\CONS/n537 ), .A(\CONS/n637 ), .B(
        \CONS/n639 ), .S(\pk_saseo_h[1] ) );
    snl_invx05 \REG_2/U127  ( .ZN(\REG_2/n410 ), .A(n10734) );
    snl_and03x1 \CODEIF/U220  ( .Z(\pgfdout[1] ), .A(\CODEIF/fm_config[1] ), 
        .B(\CODEIF/n3863 ), .C(mem_cnfg_h) );
    snl_sffqenrnx1 \LDCHK/pglpinff_reg[3]  ( .Q(\LDCHK/pglpinff[3] ), .D(1'b0), 
        .EN(1'b1), .RN(n10733), .SD(\LDCHK/lpex[3] ), .SE(ph_lpdilth), .CP(
        SCLK) );
    snl_invx05 \LBUS/U616  ( .ZN(\LBUS/n1441 ), .A(ph_lbwrh) );
    snl_and23x0 \LBUS/U631  ( .Z(\LBUS/n1436 ), .A(ph_ovfihbh), .B(
        \LBUS/n1599 ), .C(\LBUS/n1597 ) );
    snl_nand03x0 \CONS/U146  ( .ZN(\CONS/n710 ), .A(\CONS/n711 ), .B(
        \CONS/n712 ), .C(\CONS/n713 ) );
    snl_invx05 \PDOSEL/U95  ( .ZN(\PDOSEL/n105 ), .A(CDIN[51]) );
    snl_nand03x0 \CONS/U161  ( .ZN(\CONS/n746 ), .A(\CONS/n747 ), .B(
        \CONS/n748 ), .C(\CONS/n749 ) );
    snl_ffqx1 \MAIN/EXCEP_2H_reg  ( .Q(\MAIN/EXCEP_2H ), .D(\MAIN/EXCEP_1H ), 
        .CP(SCLK) );
    snl_xnor2x0 \LDCHK/U109  ( .ZN(\LDCHK/n3286 ), .A(\pgmuxout[9] ), .B(
        \pgmuxout[11] ) );
    snl_sffqenrnx1 \LBUS/ph_selldh_reg  ( .Q(ph_selldh), .D(1'b0), .EN(1'b1), 
        .RN(n10734), .SD(\pgsadrh[1] ), .SE(\LBUS/*cell*3982/U188/CONTROL1 ), 
        .CP(SCLK) );
    snl_xnor2x0 \CONS/U251  ( .ZN(\CONS/n729 ), .A(\pk_idcx_h[2] ), .B(
        \pk_indx_h[2] ) );
    snl_oai2222x0 \REGF/U368  ( .ZN(\REGF/RI_SRA12M[1] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8147 ), .C(\REGF/n8145 ), .D(\REGF/n8051 ), .E(\REGF/n8229 ), 
        .F(\REGF/n8205 ), .G(\REGF/n8230 ), .H(\REGF/n8206 ) );
    snl_oai222x0 \REGF/U439  ( .ZN(\REGF/RI_EACC[26] ), .A(\REGF/n8070 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8071 ), .E(\REGF/n8072 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U457  ( .ZN(\REGF/RI_EACC[8] ), .A(\REGF/n8124 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8125 ), .E(\REGF/n8126 ), 
        .F(\REGF/n8059 ) );
    snl_aob1b12x0 \REGF/U557  ( .Z(\REGF/RI_SRDA[0] ), .A(\REGF/n8210 ), .B(
        \pgldi[0] ), .C(\REGF/n8213 ), .D(\REGF/n8214 ) );
    snl_oai022x1 \REGF/U640  ( .ZN(\REGF/RI_TBAI[17] ), .A(\REGF/n8225 ), .B(
        \REGF/n8087 ), .C(\REGF/n8226 ), .D(\REGF/n8165 ) );
    snl_nand02x1 \ALUIS/U45  ( .ZN(\pgaluina[29] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3687 ) );
    snl_and02x1 \UPIF/U17  ( .Z(\ph_pdis_h[5] ), .A(\pk_rread_h[46] ), .B(
        \UPIF/n1046 ) );
    snl_invx05 \REGF/U667  ( .ZN(\REGF/n8120 ), .A(PDLIN[10]) );
    snl_xor2x0 \CONS/U48  ( .Z(\CONS/n570 ), .A(\pk_saco_lh[9] ), .B(
        \pgsdprlh[9] ) );
    snl_aoi022x1 \MAIN/U134  ( .ZN(\MAIN/n3621 ), .A(rmw21), .B(
        \MAIN/ph_rdwr1selh ), .C(rmw22), .D(\MAIN/ph_rdwr2selh ) );
    snl_and02x1 \UPIF/U9  ( .Z(\ph_pdis_h[4] ), .A(\pk_rread_h[55] ), .B(
        \UPIF/n1046 ) );
    snl_oai012x1 \PDOSEL/U39  ( .ZN(PDH[55]), .A(\PDOSEL/n109 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_ffqx1 \LBUS/ph_sdirlth_reg  ( .Q(ph_sdirlth), .D(ph_lbussth), .CP(SCLK
        ) );
    snl_nand04x0 \REGF/U825  ( .ZN(\REGF/n8238 ), .A(\REGF/RO_ACC[29] ), .B(
        \REGF/RO_ACC[28] ), .C(\REGF/RO_ACC[15] ), .D(\REGF/RO_ACC[19] ) );
    snl_nand02x1 \ADOSEL/U104  ( .ZN(\ADOSEL/n4140 ), .A(\pgbluext[1] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \ALUIS/U62  ( .ZN(\pgaluinb[14] ), .A(\ALUIS/n3718 ), .B(
        \ALUIS/n3719 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[4]  ( .Q(\ph_segset_h[4] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[4]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_xor2x0 \CODEIF/U297  ( .Z(\CODEIF/n3923 ), .A(\CODEIF/n3961 ), .B(
        \CODEIF/n3959 ) );
    snl_xor2x0 \CODEIF/U307  ( .Z(\CODEIF/n3977 ), .A(CDIN[30]), .B(CDIN[32])
         );
    snl_xor2x0 \CODEIF/U320  ( .Z(\CODEIF/n3997 ), .A(CDOUT[49]), .B(CDOUT[52]
        ) );
    snl_nand02x1 \ALUIS/U79  ( .ZN(\pgaluinb[31] ), .A(\ALUIS/n3752 ), .B(
        \ALUIS/n3753 ) );
    snl_aoi012x1 \ALUIS/U110  ( .ZN(\ALUIS/n3739 ), .A(\pgldi[24] ), .B(
        srcbsel), .C(allfbsel) );
    snl_nand03x0 \BLU/U357  ( .ZN(\BLU/n1533 ), .A(\BLU/n1495 ), .B(
        \BLU/n1498 ), .C(\BLU/n1492 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[10]  ( .Q(CA[10]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3851 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_invx05 \LDIS/U146  ( .ZN(\LDIS/n3125 ), .A(\pgld32[25] ) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[5]  ( .Q(\REG_2/RETCNT[5] ), .D(
        \REG_2/ph_retcnt_h[5] ), .EN(\REG_2/n517 ), .RN(\REG_2/n435 ), .SD(
        \REG_2/ncnt2[2] ), .SE(ph_d53lth), .CP(SCLK) );
    snl_oai012x1 \PDOSEL/U22  ( .ZN(PDH[38]), .A(\PDOSEL/n82 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_invx05 \LDIS/U161  ( .ZN(\LDIS/n3117 ), .A(\pgld32[17] ) );
    snl_mux21x1 \ALUSHT/U35  ( .Z(\pkdptout[17] ), .A(\ALUSHT/pkshtout[17] ), 
        .B(\ALUSHT/pkaluout[17] ), .S(\ALUSHT/n3112 ) );
    snl_oai012x1 \LBUS/U686  ( .ZN(\LBUS/n1403 ), .A(\LBUS/n1435 ), .B(
        \LBUS/n1598 ), .C(\LBUS/n1454 ) );
    snl_xor2x0 \CONS/U74  ( .Z(\CONS/n592 ), .A(\pk_pc_h[6] ), .B(
        \pk_pcs1_h[6] ) );
    snl_oai022x1 \SAEXE/U111  ( .ZN(ph_word32h), .A(\SAEXE/n413 ), .B(
        \SAEXE/n418 ), .C(\SAEXE/wrd_datah ), .D(\SAEXE/n415 ) );
    snl_mux21x1 \ALUSHT/U12  ( .Z(\pkdptout[9] ), .A(\ALUSHT/pkshtout[9] ), 
        .B(\ALUSHT/pkaluout[9] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U53  ( .Z(\CONS/n575 ), .A(\pk_saco_lh[3] ), .B(
        \pgsdprlh[3] ) );
    snl_nand02x1 \SAEXE/U136  ( .ZN(\SAEXE/n431 ), .A(\pk_psae_h[5] ), .B(
        \SAEXE/singlen ) );
    snl_aoi022x1 \ALUIS/U137  ( .ZN(\ALUIS/n3714 ), .A(\stream4[12] ), .B(
        immbsel), .C(\pk_adb_h[12] ), .D(po_brsel_h) );
    snl_nand02x1 \BLU/U370  ( .ZN(\BLU/n1489 ), .A(\BLU/n1569 ), .B(
        \BLU/n1565 ) );
    snl_xnor2x0 \LDCHK/U112  ( .ZN(\LDCHK/n3289 ), .A(\pgmuxout[13] ), .B(
        \pgmuxout[8] ) );
    snl_and02x1 \LBUS/U591  ( .Z(ph_lbe2_h), .A(phsaerrh), .B(\LBUS/OBMSEL )
         );
    snl_oai222x0 \REGF/U470  ( .ZN(\REGF/RI_DPR[23] ), .A(\REGF/n8159 ), .B(
        \REGF/n8160 ), .C(\REGF/n8161 ), .D(\REGF/n8162 ), .E(\REGF/n8081 ), 
        .F(\REGF/n8151 ) );
    snl_invx05 \REGF/U740  ( .ZN(\REGF/n8088 ), .A(\pgldi[20] ) );
    snl_invx05 \REGF/U767  ( .ZN(\REGF/n8206 ), .A(\pgsdprlh[1] ) );
    snl_nand02x1 \ADOSEL/U60  ( .ZN(\ADOSEL/n4157 ), .A(\pgsadrh[1] ), .B(
        ph_word32_h) );
    snl_ffqrnx1 \MAIN/dprw_tap1_reg  ( .Q(\MAIN/dprw_tap1 ), .D(
        \pk_rwrit_h[66] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \REGF/U802  ( .ZN(\REGF/n8089 ), .A(\pkdptout[20] ) );
    snl_invx05 \ADOSEL/U47  ( .ZN(\ADOSEL/n4117 ), .A(\pkdptout[9] ) );
    snl_and02x1 \LDCHK/U96  ( .Z(\LDCHK/n3274 ), .A(ph_word32_h), .B(
        \pgsadrh[0] ) );
    snl_or02x1 \PDOSEL/U151  ( .Z(\PDOSEL/n226 ), .A(mem_cnfg_h), .B(
        write_pr_h) );
    snl_ffqrnx1 \LBUS/phsaerrh_reg  ( .Q(phsaerrh), .D(ph_lberr), .RN(n10734), 
        .CP(SCLK) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[3]  ( .Q(\CODEIF/pfctr[3] ), .D(
        \CODEIF/pfctr415[3] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_oai112x0 \LBUS/U644  ( .ZN(\LBUS/n1422 ), .A(ph_ovfihbh), .B(
        \LBUS/n1599 ), .C(\LBUS/n1435 ), .D(\LBUS/n1597 ) );
    snl_nor03x0 \CONS/U133  ( .ZN(\CONS/n674 ), .A(\CONS/n588 ), .B(
        \CONS/n586 ), .C(\CONS/n587 ) );
    snl_oai122x0 \ADOSEL/U29  ( .ZN(\pgmuxout[18] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4096 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4095 ), .E(
        \ADOSEL/n4141 ) );
    snl_invx05 \CODEIF/U272  ( .ZN(\CODEIF/n3920 ), .A(\CODEIF/pfctr[18] ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[10]  ( .Q(\CODEIF/pfctr[10] ), .D(
        \CODEIF/pfctr415[10] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_muxi21x1 \LDIS/U184  ( .ZN(\LDIS/ldexch[26] ), .A(\LDIS/n3162 ), .B(
        \LDIS/n3161 ), .S(\LDIS/n3165 ) );
    snl_oai013x0 \LBUS/U574  ( .ZN(\LBUS/nlt[3] ), .A(\LBUS/n1416 ), .B(
        ph_timouth), .C(LDS), .D(\LBUS/n1430 ) );
    snl_xnor2x0 \CONS/U203  ( .ZN(\CONS/n690 ), .A(\pk_pc_h[7] ), .B(
        \pk_pcs2_h[7] ) );
    snl_and02x1 \REG_2/U152  ( .Z(\ph_cpudout[22] ), .A(\ph_segset_h[22] ), 
        .B(seg_cnfg_h) );
    snl_nand02x1 \BLU/U395  ( .ZN(\BLU/n1474 ), .A(\BLU/n1567 ), .B(
        \BLU/n1563 ) );
    snl_oa2222x1 \BLU/U414  ( .Z(\BLU/n1515 ), .A(\BLU/n1498 ), .B(\BLU/n1500 
        ), .C(\BLU/n1495 ), .D(\BLU/n1497 ), .E(\BLU/n1492 ), .F(\BLU/n1494 ), 
        .G(\BLU/n1489 ), .H(\BLU/n1491 ) );
    snl_oai222x0 \REGF/U445  ( .ZN(\REGF/RI_EACC[20] ), .A(\REGF/n8088 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8089 ), .E(\REGF/n8090 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U487  ( .ZN(\REGF/RI_DPR[6] ), .A(\REGF/n8195 ), .B(
        \REGF/n8160 ), .C(\REGF/n8196 ), .D(\REGF/n8162 ), .E(\REGF/n8132 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U495  ( .Z(\REGF/RI_PCOL[30] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[30]), .C(\stream4[30] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U635  ( .Z(\REGF/RI_STAT[0] ), .A(PDLIN[0]), .B(
        \ph_pdis_h[4] ), .C(obacc), .D(\REGF/n8224 ) );
    snl_invx05 \REGF/U699  ( .ZN(\REGF/n8099 ), .A(PDLIN[17]) );
    snl_nand02x1 \CODEIF/U255  ( .ZN(\CODEIF/n3867 ), .A(cnt_write_h), .B(
        \CODEIF/n3944 ) );
    snl_oa023x1 \LBUS/U553  ( .Z(\LBUS/n1392 ), .A(\LBUS/n1419 ), .B(
        \LBUS/ilt[0] ), .C(\LBUS/n1420 ), .D(\LBUS/n1421 ), .E(\LBUS/n1422 )
         );
    snl_xnor2x0 \CONS/U224  ( .ZN(\CONS/n713 ), .A(\pk_idcz_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_invx05 \BLU/U433  ( .ZN(\BLU/n1527 ), .A(allfbsel) );
    snl_invx05 \LBUS/U663  ( .ZN(\LBUS/n1406 ), .A(\LBUS/n1435 ) );
    snl_xor2x0 \CONS/U91  ( .Z(\CONS/n609 ), .A(\pk_idcz_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_invx05 \REGF/U709  ( .ZN(\REGF/n8223 ), .A(\ph_pdis_h[4] ) );
    snl_ao022x1 \MAIN/U166  ( .Z(\MAIN/n3633 ), .A(\MAIN/ph_rdwr2selh ), .B(
        saenabl2), .C(\MAIN/ph_rdwr1selh ), .D(saenabl1) );
    snl_xor2x0 \CONS/U114  ( .Z(\CONS/n632 ), .A(\pk_idcw_h[15] ), .B(
        \pk_indw_h[15] ) );
    snl_nor02x1 \PDOSEL/U118  ( .ZN(\PDOSEL/n149 ), .A(\ph_cpudout[24] ), .B(
        \pk_pdo_h[24] ) );
    snl_nand02x1 \CODEIF/U369  ( .ZN(\CODEIF/n3963 ), .A(\CODEIF/fm_config[0] 
        ), .B(\CODEIF/n3863 ) );
    snl_invx1 \ALUIS/U30  ( .ZN(\ALUIS/n3657 ), .A(allfasel) );
    snl_nand02x1 \ALUIS/U159  ( .ZN(\ALUIS/n3682 ), .A(\pk_ada_h[24] ), .B(
        po_arsel_h) );
    snl_xor2x0 \LDCHK/U73  ( .Z(\LDCHK/n3302 ), .A(\pgld32[22] ), .B(
        \pgld32[21] ) );
    snl_ao022x1 \REGF/U505  ( .Z(\REGF/RI_PCOL[20] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[20]), .C(\stream4[20] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U517  ( .Z(\REGF/RI_PCOL[8] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[8]), .C(\stream4[8] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U522  ( .Z(\REGF/RI_PCOL[3] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[3]), .C(\stream4[3] ), .D(\REGF/n8209 ) );
    snl_invx1 \ALUIS/U17  ( .ZN(\pgaluina[14] ), .A(\ALUIS/n3649 ) );
    snl_ffqrnx1 \MAIN/sprw_tap2_reg  ( .Q(\MAIN/sprw_tap2 ), .D(
        \MAIN/sprw_tap1 ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \LDIS/U218  ( .ZN(\LDIS/n3160 ), .A(LIN[27]) );
    snl_aoi122x0 \BLU/U339  ( .ZN(\BLU/n1524 ), .A(\pk_stat_h[0] ), .B(accbsel
        ), .C(pk_bitdatah), .D(srcbsel), .E(\BLU/n1554 ) );
    snl_oai222x0 \REGF/U612  ( .ZN(\REGF/RI_SPR[17] ), .A(\REGF/n8173 ), .B(
        \REGF/n8220 ), .C(\REGF/n8174 ), .D(\REGF/n8221 ), .E(\REGF/n8099 ), 
        .F(\REGF/n8218 ) );
    snl_nand02x1 \ADOSEL/U85  ( .ZN(\ADOSEL/n4106 ), .A(\pgbluext[5] ), .B(
        \ADOSEL/n4156 ) );
    snl_oai012x1 \LDIS/U128  ( .ZN(\pgldi[15] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3114 ), .C(\LDIS/n3115 ) );
    snl_or02x1 \MAIN/U141  ( .Z(\MAIN/cstregw_inhibith ), .A(
        \MAIN/cstregw_tap2 ), .B(\MAIN/cstregw_tap1 ) );
    snl_muxi21x1 \LDCHK/U54  ( .ZN(\LDCHK/lpex[1] ), .A(\LDCHK/n3273 ), .B(
        \LDCHK/n3272 ), .S(\LDCHK/n3277 ) );
    snl_oai222x0 \REGF/U627  ( .ZN(\REGF/RI_SPR[2] ), .A(\REGF/n8203 ), .B(
        \REGF/n8220 ), .C(\REGF/n8204 ), .D(\REGF/n8221 ), .E(\REGF/n8144 ), 
        .F(\REGF/n8218 ) );
    snl_and12x1 \REGF/U782  ( .Z(\REGF/n8053 ), .A(\ph_pdis_h[5] ), .B(
        ph_rgfile_h) );
    snl_xor2x0 \LDCHK/U61  ( .Z(\LDCHK/n3261 ), .A(\LDCHK/n3288 ), .B(
        \LDCHK/n3289 ) );
    snl_invx05 \PDOSEL/U79  ( .ZN(\PDOSEL/n94 ), .A(CDIN[40]) );
    snl_nand02x2 \ALUIS/U22  ( .ZN(\pgaluina[13] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3671 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[0]  ( .Q(\ph_segset_h[0] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[0]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_ao2222x1 \REGF/U530  ( .Z(\REGF/RI_SRDA[27] ), .A(PDLIN[27]), .B(
        \ph_pdis_h[9] ), .C(\pgldi[27] ), .D(\REGF/n8210 ), .E(\stream3[27] ), 
        .F(\REGF/n8211 ), .G(\pkdptout[27] ), .H(\REGF/n8212 ) );
    snl_sffqenrnx1 \LBUS/PIOSEL_1_reg  ( .Q(\LBUS/PIOSEL_1_Q1249 ), .D(1'b0), 
        .EN(1'b1), .RN(n10734), .SD(\LBUS/*cell*3982/U31/CONTROL1 ), .SE(
        \LBUS/*cell*3982/U185/CONTROL1 ), .CP(SCLK) );
    snl_oai222x0 \REGF/U600  ( .ZN(\REGF/RI_ACC[1] ), .A(\REGF/n8145 ), .B(
        \REGF/n8215 ), .C(\REGF/n8146 ), .D(\REGF/n8216 ), .E(\REGF/n8147 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U790  ( .ZN(\REGF/n8057 ), .A(\pkdptout[31] ) );
    snl_nand02x1 \ADOSEL/U97  ( .ZN(\ADOSEL/n4146 ), .A(\pgbluext[7] ), .B(
        \ADOSEL/n4156 ) );
    snl_aoi012x1 \MAIN/U153  ( .ZN(\MAIN/n3622 ), .A(\MAIN/n3634 ), .B(
        \MAIN/n3632 ), .C(\MAIN/ph_rrmwh ) );
    snl_xor2x0 \CODEIF/U247  ( .Z(CPOUT[1]), .A(\CODEIF/n3940 ), .B(
        \CODEIF/n3941 ) );
    snl_invx05 \CODEIF/U260  ( .ZN(\CODEIF/n3884 ), .A(\CODEIF/pfctr[6] ) );
    snl_xor2x0 \LDCHK/U46  ( .Z(\LDCHK/n3233 ), .A(\LDCHK/n3260 ), .B(
        \LDCHK/n3261 ) );
    snl_invx05 \LDIS/U196  ( .ZN(\LDIS/n3164 ), .A(LIN[16]) );
    snl_invx05 \LBUS/U656  ( .ZN(\LBUS/n1593 ), .A(\LBUS/n1462 ) );
    snl_nor02x1 \LBUS/U566  ( .ZN(ph_pdhen_h), .A(\LBUS/n1411 ), .B(
        \LBUS/n1391 ) );
    snl_aoi023x0 \CONS/U121  ( .ZN(\CONS/n641 ), .A(\CONS/n642 ), .B(
        \CONS/n643 ), .C(\CONS/n644 ), .D(\CONS/n645 ), .E(\CONS/n646 ) );
    snl_invx05 \BLU/U387  ( .ZN(\BLU/n1467 ), .A(\pgld16[15] ) );
    snl_xnor2x0 \CONS/U211  ( .ZN(\CONS/n694 ), .A(\pk_pc_h[7] ), .B(
        \pk_pcs1_h[7] ) );
    snl_and02x1 \REG_2/U140  ( .Z(\ph_cpudout[10] ), .A(\ph_segset_h[10] ), 
        .B(seg_cnfg_h) );
    snl_aoi112x0 \BLU/U406  ( .ZN(\BLU/n1577 ), .A(\poalufnc[0] ), .B(
        \BLU/n1552 ), .C(\BLU/n1525 ), .D(\poalufnc[1] ) );
    snl_nand04x0 \LBUS/U671  ( .ZN(\LBUS/n1432 ), .A(LBER), .B(\LBUS/n1601 ), 
        .C(\LBUS/temp[3] ), .D(\LBUS/n1459 ) );
    snl_xor2x0 \CONS/U83  ( .Z(\CONS/n601 ), .A(\pk_idcz_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_xnor2x0 \CONS/U236  ( .ZN(\CONS/n717 ), .A(\pk_idcy_h[17] ), .B(
        \pk_indy_h[17] ) );
    snl_invx05 \BLU/U421  ( .ZN(\BLU/n1537 ), .A(\BLU/n1492 ) );
    snl_xor2x0 \CONS/U106  ( .Z(\CONS/n624 ), .A(\pk_idcx_h[13] ), .B(
        \pk_indx_h[13] ) );
    snl_oai222x0 \REGF/U462  ( .ZN(\REGF/RI_EACC[3] ), .A(\REGF/n8139 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8140 ), .E(\REGF/n8141 ), 
        .F(\REGF/n8059 ) );
    snl_invx05 \REGF/U752  ( .ZN(\REGF/n8148 ), .A(\pgldi[0] ) );
    snl_invx05 \REGF/U775  ( .ZN(\REGF/n8182 ), .A(\pgsdprlh[13] ) );
    snl_oai122x0 \CODEIF/U229  ( .ZN(\CODEIF/pfctr415[8] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3890 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3891 ), .E(
        \CODEIF/n3892 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[1]  ( .Q(CA[1]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3842 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_xnor2x0 \CONS/U258  ( .ZN(\CONS/n347 ), .A(\pk_idcx_h[0] ), .B(
        \pk_indx_h[0] ) );
    snl_invx05 \ADOSEL/U72  ( .ZN(\ADOSEL/n4125 ), .A(\pkdptout[28] ) );
    snl_xnor2x0 \CONS/U168  ( .ZN(\CONS/n556 ), .A(\pk_saco_hh[30] ), .B(
        \pgsdprhh[30] ) );
    snl_nor04x0 \LDCHK/U84  ( .ZN(\LDCHK/n3242 ), .A(\pgld32[7] ), .B(
        \pgld32[4] ), .C(\pgld32[13] ), .D(\pgld32[2] ) );
    snl_oa012x1 \LBUS/U638  ( .Z(\LBUS/n1428 ), .A(\LBUS/ilt[0] ), .B(
        \LBUS/n1453 ), .C(\LBUS/n1446 ) );
    snl_aoi022x1 \PDOSEL/U164  ( .ZN(\PDOSEL/n224 ), .A(PA02), .B(SWIT_wire), 
        .C(\PDOSEL/n225 ), .D(\PDOSEL/n76 ) );
    snl_invx05 \ADOSEL/U55  ( .ZN(\ADOSEL/n4105 ), .A(\pkdptout[5] ) );
    snl_nand02x1 \PDOSEL/U143  ( .ZN(\PDOSEL/n134 ), .A(CDIN[27]), .B(
        \PDOSEL/n119 ) );
    snl_oai022x1 \REGF/U649  ( .ZN(\REGF/RI_TBAI[5] ), .A(\REGF/n8225 ), .B(
        \REGF/n8123 ), .C(\REGF/n8226 ), .D(\REGF/n8189 ) );
    snl_invx05 \REGF/U810  ( .ZN(\REGF/n8110 ), .A(\pkdptout[13] ) );
    snl_ffqsnx1 \CODEIF/pgfddacntl_reg  ( .Q(CDCNT), .D(\CODEIF/fddacnt_in ), 
        .SN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_xor2x0 \CODEIF/U332  ( .Z(\CODEIF/n4013 ), .A(CDOUT[21]), .B(CDOUT[19]
        ) );
    snl_aoi012x1 \ALUIS/U102  ( .ZN(\ALUIS/n3747 ), .A(\pgldi[28] ), .B(
        srcbsel), .C(allfbsel) );
    snl_invx05 \BLU/U345  ( .ZN(\BLU/n1560 ), .A(\pgbitnoh[1] ) );
    snl_invx05 \LDIS/U154  ( .ZN(\LDIS/n3114 ), .A(\pgld32[15] ) );
    snl_muxi21x1 \LDIS/U173  ( .ZN(\LDIS/ldexcl[14] ), .A(\LDIS/n3153 ), .B(
        \LDIS/n3154 ), .S(\LDIS/n3134 ) );
    snl_mux21x1 \ALUSHT/U27  ( .Z(\pkdptout[24] ), .A(\ALUSHT/pkshtout[24] ), 
        .B(\ALUSHT/pkaluout[24] ), .S(\ALUSHT/n3112 ) );
    snl_aoi022x1 \LBUS/U694  ( .ZN(\LBUS/n1611 ), .A(\LBUS/word32odphase ), 
        .B(\pgsadrh[1] ), .C(\LBUS/n1609 ), .D(\LBUS/n1632 ) );
    snl_xor2x0 \CONS/U66  ( .Z(\CONS/n583 ), .A(\CONS/SACO[3] ), .B(
        \pgsdprlh[7] ) );
    snl_oai012x1 \PDOSEL/U30  ( .ZN(PDH[46]), .A(\PDOSEL/n100 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nor02x1 \SAEXE/U103  ( .ZN(\SAEXE/n412 ), .A(\SAEXE/trsc2_h ), .B(
        \SAEXE/trsc1_h ) );
    snl_oai012x1 \PDOSEL/U17  ( .ZN(PDH[33]), .A(\PDOSEL/n77 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_invx05 \SAEXE/U124  ( .ZN(\SAEXE/n423 ), .A(\SAEXE/stage_2nd ) );
    snl_invx05 \CODEIF/U285  ( .ZN(\CODEIF/n3903 ), .A(PDLIN[12]) );
    snl_invx05 \CONS/U41  ( .ZN(\CONS/n546 ), .A(\pk_saco_lh[4] ) );
    snl_invx05 \BLU/U362  ( .ZN(\BLU/n1485 ), .A(\pgld16[9] ) );
    snl_xor2x0 \CODEIF/U315  ( .Z(\CODEIF/n3989 ), .A(\CODEIF/n3990 ), .B(
        \CODEIF/n3991 ) );
    snl_aoi022x1 \ALUIS/U125  ( .ZN(\ALUIS/n3726 ), .A(\stream4[18] ), .B(
        immbsel), .C(\pk_adb_h[18] ), .D(po_brsel_h) );
    snl_nand02x1 \LDCHK/U100  ( .ZN(\LDCHK/n3271 ), .A(\pgld32[29] ), .B(
        \LDCHK/n3255 ) );
    snl_invx05 \LBUS/U583  ( .ZN(\LBUS/n1632 ), .A(\pgsadrh[1] ) );
    snl_oai022x1 \REGF/U373  ( .ZN(\REGF/RI_TBAI[10] ), .A(\REGF/n8225 ), .B(
        \REGF/n8108 ), .C(\REGF/n8226 ), .D(\REGF/n8179 ) );
    snl_oai222x0 \REGF/U579  ( .ZN(\REGF/RI_ACC[22] ), .A(\REGF/n8082 ), .B(
        \REGF/n8215 ), .C(\REGF/n8083 ), .D(\REGF/n8216 ), .E(\REGF/n8084 ), 
        .F(\REGF/n8217 ) );
    snl_ao2222x1 \REGF/U545  ( .Z(\REGF/RI_SRDA[12] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[12]), .C(\pgldi[12] ), .D(\REGF/n8210 ), .E(\stream3[12] ), .F(
        \REGF/n8211 ), .G(\pkdptout[12] ), .H(\REGF/n8212 ) );
    snl_and02x1 \REGF/U562  ( .Z(\REGF/RO_LPSAS2156[4] ), .A(ph_sastlth), .B(
        \REGF/RO_EST1[6] ) );
    snl_oai022x1 \REGF/U652  ( .ZN(\REGF/RI_TBAI[2] ), .A(\REGF/n8225 ), .B(
        \REGF/n8132 ), .C(\REGF/n8226 ), .D(\REGF/n8195 ) );
    snl_nand02x1 \ALUIS/U57  ( .ZN(\pgaluinb[9] ), .A(\ALUIS/n3708 ), .B(
        \ALUIS/n3709 ) );
    snl_aoi012x1 \LBUS/U598  ( .ZN(\LBUS/n1451 ), .A(ph_lbussth), .B(
        \LBUS/ilt[4] ), .C(pgfbadrsel) );
    snl_invx05 \BLU/U379  ( .ZN(\BLU/n1503 ), .A(\pgld16[3] ) );
    snl_invx05 \REGF/U675  ( .ZN(\REGF/n8132 ), .A(PDLIN[6]) );
    snl_nor02x1 \LDCHK/U33  ( .ZN(LPOUT[2]), .A(\LDCHK/n3231 ), .B(
        \LDCHK/n3234 ) );
    snl_muxi21x1 \LDIS/U168  ( .ZN(\LDIS/ldexcl[4] ), .A(\LDIS/n3143 ), .B(
        \LDIS/n3144 ), .S(\LDIS/n3134 ) );
    snl_nor04x0 \SAEXE/U118  ( .ZN(ph_sprsel2_h), .A(\SAEXE/n427 ), .B(
        \SAEXE/n413 ), .C(\SAEXE/n428 ), .D(\SAEXE/n422 ) );
    snl_nand02x1 \MAIN/U126  ( .ZN(\MAIN/*cell*4603/U16/CONTROL1 ), .A(
        \MAIN/n3616 ), .B(\MAIN/n3617 ) );
    snl_ao022x1 \REGF/U430  ( .Z(\REGF/RI_PCOH[3] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[3]), .C(\stream4[35] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U479  ( .ZN(\REGF/RI_DPR[14] ), .A(\REGF/n8179 ), .B(
        \REGF/n8160 ), .C(\REGF/n8180 ), .D(\REGF/n8162 ), .E(\REGF/n8108 ), 
        .F(\REGF/n8151 ) );
    snl_aoi022x4 \CODEIF/U215  ( .ZN(\CODEIF/n3864 ), .A(\CODEIF/n3944 ), .B(
        \CODEIF/n4030 ), .C(\CODEIF/wpfcinc ), .D(cnt_write_h) );
    snl_xor2x0 \CODEIF/U329  ( .Z(\CODEIF/n4008 ), .A(\CODEIF/n4009 ), .B(
        \CODEIF/n4010 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[8]  ( .Q(CA[8]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3849 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_aoi022x1 \ALUIS/U119  ( .ZN(\ALUIS/n3730 ), .A(\stream4[20] ), .B(
        immbsel), .C(\pk_adb_h[20] ), .D(po_brsel_h) );
    snl_nand02x1 \ALUIS/U70  ( .ZN(\pgaluinb[22] ), .A(\ALUIS/n3734 ), .B(
        \ALUIS/n3735 ) );
    snl_xnor2x0 \CONS/U264  ( .ZN(\CONS/n740 ), .A(\pk_idcw_h[9] ), .B(
        \pk_indw_h[9] ) );
    snl_ao022x1 \REG_2/U135  ( .Z(\ph_cpudout[5] ), .A(\ph_segset_h[5] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[5] ), .D(ret_cont_h) );
    snl_xnor2x0 \CODEIF/U385  ( .ZN(\CODEIF/n3980 ), .A(CDIN[28]), .B(CDIN[29]
        ) );
    snl_xor2x0 \CODEIF/U404  ( .Z(\CODEIF/n4023 ), .A(\CODEIF/n4037 ), .B(
        CDOUT[54]) );
    snl_sffqenrnx1 \CODEIF/fm_config_reg[0]  ( .Q(\CODEIF/fm_config[0] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEIF/n3862 ), .SD(PDLIN[0]), .SE(cnfg_write_h
        ), .CP(SCLK) );
    snl_invx05 \REGF/U690  ( .ZN(\REGF/n8165 ), .A(\pgregadrh[21] ) );
    snl_invx05 \REGF/U700  ( .ZN(\REGF/n8175 ), .A(\pgregadrh[16] ) );
    snl_invx05 \REGF/U749  ( .ZN(\REGF/n8112 ), .A(\pgldi[12] ) );
    snl_nor03x0 \CONS/U154  ( .ZN(\CONS/n349 ), .A(\CONS/n624 ), .B(
        \CONS/n622 ), .C(\CONS/n623 ) );
    snl_nand02x1 \PDOSEL/U158  ( .ZN(\PDOSEL/n142 ), .A(CDIN[14]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \PDOSEL/U87  ( .ZN(\PDOSEL/n112 ), .A(CDIN[58]) );
    snl_invx05 \ADOSEL/U69  ( .ZN(\ADOSEL/n4129 ), .A(\pkdptout[13] ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[14]  ( .Q(\CODEIF/pfctr[14] ), .D(
        \CODEIF/pfctr415[14] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_invx05 \LBUS/U623  ( .ZN(\LBUS/n1415 ), .A(ph_timouth) );
    snl_oai122x0 \CODEIF/U232  ( .ZN(\CODEIF/pfctr415[11] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3899 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3900 ), .E(
        \CODEIF/n3901 ) );
    snl_xor2x0 \CODEIF/U423  ( .Z(\CODEIF/n4044 ), .A(\CODEIF/n4019 ), .B(
        \CODEIF/n4015 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[7]  ( .Q(\CODEIF/pfctr[7] ), .D(
        \CODEIF/pfctr415[7] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nor02x1 \LBUS/U604  ( .ZN(\LBUS/n1457 ), .A(ph_bit_h), .B(ph_word16_h)
         );
    snl_xnor2x0 \CONS/U173  ( .ZN(\CONS/n651 ), .A(\pgsdprlh[22] ), .B(
        \pk_saco_lh[22] ) );
    snl_xnor2x0 \CONS/U243  ( .ZN(\CONS/n521 ), .A(\pk_idcy_h[0] ), .B(
        \pk_indy_h[0] ) );
    snl_xor2x0 \CONS/U98  ( .Z(\CONS/n616 ), .A(\pk_idcy_h[14] ), .B(
        \pk_indy_h[14] ) );
    snl_nor02x1 \PDOSEL/U111  ( .ZN(\PDOSEL/n163 ), .A(\pk_pdo_h[5] ), .B(
        \ph_cpudout[5] ) );
    snl_aoi022x1 \ALUIS/U95  ( .ZN(\ALUIS/n3752 ), .A(\stream4[31] ), .B(
        immbsel), .C(\pk_adb_h[31] ), .D(po_brsel_h) );
    snl_oai2222x0 \REGF/U353  ( .ZN(\REGF/RI_SRA12M[22] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8084 ), .C(\REGF/n8082 ), .D(\REGF/n8051 ), .E(\REGF/n8163 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8164 ) );
    snl_oai222x2 \REGF/U391  ( .ZN(\REGF/RI_SRA12M[26] ), .A(\REGF/n8060 ), 
        .B(\REGF/n8051 ), .C(\REGF/n8227 ), .D(\REGF/n8154 ), .E(\REGF/n8228 ), 
        .F(\REGF/n8062 ) );
    snl_nand02x2 \REGF/U396  ( .ZN(\REGF/n8226 ), .A(ph_tprsel_h), .B(
        \REGF/n8225 ) );
    snl_oai222x0 \REGF/U587  ( .ZN(\REGF/RI_ACC[14] ), .A(\REGF/n8106 ), .B(
        \REGF/n8215 ), .C(\REGF/n8107 ), .D(\REGF/n8216 ), .E(\REGF/n8108 ), 
        .F(\REGF/n8217 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[9]  ( .Q(\ph_segset_h[9] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n435 ), .SD(PDLIN[9]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_ao022x1 \REGF/U410  ( .Z(\REGF/RI_PCOH[23] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[23]), .C(\stream4[55] ), .D(\REGF/n8053 ) );
    snl_ao022x1 \REGF/U417  ( .Z(\REGF/RI_PCOH[16] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[16]), .C(\stream4[48] ), .D(\REGF/n8053 ) );
    snl_invx05 \REGF/U720  ( .ZN(\REGF/n8136 ), .A(\pgldi[4] ) );
    snl_invx05 \REGF/U727  ( .ZN(\REGF/n8063 ), .A(\pgldi[29] ) );
    snl_oai122x0 \ADOSEL/U20  ( .ZN(\pgmuxout[9] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4116 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4117 ), .E(
        \ADOSEL/n4118 ) );
    snl_ffqrnx1 \LBUS/ph_lbusylth_reg  ( .Q(\LBUS/ph_lbusylth ), .D(LBSY), 
        .RN(n10734), .CP(SCLK) );
    snl_nand02x1 \PDOSEL/U136  ( .ZN(\PDOSEL/n180 ), .A(CDIN[8]), .B(
        \PDOSEL/n119 ) );
    snl_nand02x1 \CODEIF/U347  ( .ZN(\CODEIF/n3871 ), .A(\CODEIF/pgctrinc[1] ), 
        .B(\CODEIF/n3945 ) );
    snl_invx05 \MAIN/U148  ( .ZN(\MAIN/n3627 ), .A(\MAIN/ph_rdwr1selh ) );
    snl_ao022x1 \LDIS/U121  ( .Z(\pgld16[11] ), .A(ph_selldl), .B(\pgld32[11] 
        ), .C(ph_selldh), .D(\pgld32[27] ) );
    snl_sffqenrnx1 \LBUS/OBMSEL_reg  ( .Q(\LBUS/OBMSEL ), .D(1'b0), .EN(1'b1), 
        .RN(n10734), .SD(ph_obmselh), .SE(\LBUS/n1393 ), .CP(SCLK) );
    snl_invx05 \CMPX/U30  ( .ZN(ph_adrinc_h), .A(\CMPX/n1049 ) );
    snl_xnor2x0 \CONS/U196  ( .ZN(\CONS/n675 ), .A(\pk_pc_h[15] ), .B(
        \pk_pcs2_h[15] ) );
    snl_oai112x0 \PDOSEL/U45  ( .ZN(PDLOUT[25]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n111 ), .C(\PDOSEL/n117 ), .D(\PDOSEL/n118 ) );
    snl_sffqenrnx1 \LBUS/MMBSEL_reg  ( .Q(\LBUS/MMBSEL ), .D(1'b0), .EN(1'b1), 
        .RN(n10734), .SD(ph_mmbselh), .SE(\LBUS/n1393 ), .CP(SCLK) );
    snl_nor02x1 \BLU/U330  ( .ZN(\BLU/n1508 ), .A(\BLU/n1543 ), .B(\BLU/n1542 
        ) );
    snl_xor2x0 \CODEIF/U360  ( .Z(\CODEIF/n3955 ), .A(CDIN[24]), .B(
        \CODEIF/n3952 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[14]  ( .Q(CA[14]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3861 ), .SD(\CODEIF/n3855 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_invx05 \LDIS/U211  ( .ZN(\LDIS/n3135 ), .A(LIN[8]) );
    snl_nand02x1 \ALUIS/U150  ( .ZN(\ALUIS/n3661 ), .A(\pk_ada_h[3] ), .B(
        po_arsel_h) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[1]  ( .Q(\REG_2/RETCNT[1] ), .D(
        \REG_2/ph_retcnt_h[1] ), .EN(\REG_2/n517 ), .RN(\REG_2/n435 ), .SD(
        \REG_2/ncnt1[1] ), .SE(ph_d20lth), .CP(SCLK) );
    snl_nand02x1 \ALUIS/U39  ( .ZN(\pgaluina[23] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3681 ) );
    snl_ao022x1 \BLUOS/U20  ( .Z(\pgbluext[1] ), .A(\pkbludgh[1] ), .B(
        ph_bit_h), .C(\pkdptout[1] ), .D(ph_word16_h) );
    snl_aoi013x0 \CONS/U34  ( .ZN(\CONS/n539 ), .A(\pk_saco_lh[4] ), .B(
        \CONS/n540 ), .C(\CONS/n541 ), .D(\CONS/n542 ) );
    snl_nand04x0 \BLU/U317  ( .ZN(\BLU/SRC_DATA_M ), .A(\BLU/n1513 ), .B(
        \BLU/n1514 ), .C(\BLU/n1515 ), .D(\BLU/n1516 ) );
    snl_ao022x1 \LDIS/U106  ( .Z(\pgldi[4] ), .A(ph_word32_h), .B(\pgld32[4] ), 
        .C(\pgld16[4] ), .D(ph_word16_h) );
    snl_nand02x1 \CMPX/U17  ( .ZN(ph_adrwtenh), .A(\CMPX/n1049 ), .B(
        \CMPX/n1050 ) );
    snl_oai112x0 \PDOSEL/U62  ( .ZN(PDLOUT[24]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n110 ), .C(\PDOSEL/n148 ), .D(\PDOSEL/n149 ) );
    snl_oai122x0 \ADOSEL/U27  ( .ZN(\pgmuxout[16] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4090 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4088 ), .E(
        \ADOSEL/n4139 ) );
    snl_nor02x1 \PDOSEL/U131  ( .ZN(\PDOSEL/n137 ), .A(\ph_cpudout[12] ), .B(
        \pk_pdo_h[12] ) );
    snl_ao2b2b2x0 \REGF/U437  ( .Z(\REGF/RI_EACC[28] ), .A(\REGF/n8065 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8066 ), .E(PDLIN[28]), .F(
        \ph_pdis_h[1] ) );
    snl_oai222x0 \REGF/U580  ( .ZN(\REGF/RI_ACC[21] ), .A(\REGF/n8085 ), .B(
        \REGF/n8215 ), .C(\REGF/n8086 ), .D(\REGF/n8216 ), .E(\REGF/n8087 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U697  ( .ZN(\REGF/n8096 ), .A(PDLIN[18]) );
    snl_aoi012x1 \ALUIS/U92  ( .ZN(\ALUIS/n3697 ), .A(\pgldi[3] ), .B(srcbsel), 
        .C(allfbsel) );
    snl_invx05 \REGF/U707  ( .ZN(\REGF/n8138 ), .A(PDLIN[4]) );
    snl_nand02x1 \ADOSEL/U111  ( .ZN(\ADOSEL/n4121 ), .A(\pgbluext[26] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \CODEIF/U340  ( .ZN(\CODEIF/n3892 ), .A(\CODEIF/pgctrinc[8] ), 
        .B(\CODEIF/n3945 ) );
    snl_xor2x0 \CODEIF/U367  ( .Z(\CODEIF/n4028 ), .A(\CODEIF/n4029 ), .B(
        \CODEIF/n4020 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[16]  ( .Q(CA[16]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3857 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_ffqrnx1 \CODEIF/pgiaendp_reg  ( .Q(pgiaendp), .D(\CODEIF/friend_in ), 
        .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_ao022x1 \BLUOS/U27  ( .Z(\pgbluext[8] ), .A(\pkbludgh[8] ), .B(
        ph_bit_h), .C(\pkdptout[8] ), .D(ph_word16_h) );
    snl_invx05 \MAIN/U168  ( .ZN(\MAIN/ph_rmw1h ), .A(\MAIN/n3620 ) );
    snl_oai112x0 \PDOSEL/U65  ( .ZN(PDLOUT[22]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n108 ), .C(\PDOSEL/n154 ), .D(\PDOSEL/n155 ) );
    snl_nor02x1 \PDOSEL/U116  ( .ZN(\PDOSEL/n141 ), .A(\ph_cpudout[26] ), .B(
        \pk_pdo_h[26] ) );
    snl_ao022x1 \LDIS/U101  ( .Z(\pgld16[1] ), .A(ph_selldl), .B(\pgld32[1] ), 
        .C(ph_selldh), .D(\pgld32[17] ) );
    snl_nand12x1 \CMPX/U10  ( .ZN(ph_locken_h), .A(ph_lockh), .B(\CMPX/n1048 )
         );
    snl_and02x1 \CONS/U33  ( .Z(ph_pccons_h), .A(\CONS/n538 ), .B(pk_pcsee_h)
         );
    snl_oai022x1 \BLU/U310  ( .ZN(\pkbludgh[6] ), .A(\BLU/n1464 ), .B(
        \BLU/n1492 ), .C(\BLU/n1493 ), .D(\BLU/n1494 ) );
    snl_and02x1 \ALUIS/U19  ( .Z(\ALUIS/n3651 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3663 ) );
    snl_nand02x1 \ALUIS/U157  ( .ZN(\ALUIS/n3684 ), .A(\pk_ada_h[26] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U216  ( .ZN(\LDIS/n3162 ), .A(LIN[26]) );
    snl_nand02x1 \ALUIS/U77  ( .ZN(\pgaluinb[29] ), .A(\ALUIS/n3748 ), .B(
        \ALUIS/n3749 ) );
    snl_nand02x1 \ALUIS/U170  ( .ZN(\ALUIS/n3672 ), .A(\pk_ada_h[14] ), .B(
        po_arsel_h) );
    snl_ao022x1 \LDIS/U126  ( .Z(\pgldi[14] ), .A(ph_word32_h), .B(
        \pgld32[14] ), .C(\pgld16[14] ), .D(ph_word16_h) );
    snl_xnor2x0 \CONS/U191  ( .ZN(\CONS/n671 ), .A(\pgsdprlh[22] ), .B(
        \CONS/SACO[18] ) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[3]  ( .Q(\REG_2/RETCNT[3] ), .D(
        \REG_2/ph_retcnt_h[3] ), .EN(\REG_2/n517 ), .RN(\REG_2/n435 ), .SD(
        \REG_2/ncnt2[0] ), .SE(ph_d53lth), .CP(SCLK) );
    snl_nor04x0 \BLU/U337  ( .ZN(\BLU/n1511 ), .A(\BLU/n1541 ), .B(\BLU/n1543 
        ), .C(\BLU/n1551 ), .D(\BLU/n1540 ) );
    snl_oai012x1 \PDOSEL/U42  ( .ZN(PDH[58]), .A(\PDOSEL/n112 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nor04x0 \BLU/U359  ( .ZN(\BLU/n1571 ), .A(\BLU/n1533 ), .B(\BLU/n1539 
        ), .C(\BLU/n1538 ), .D(\BLU/n1551 ) );
    snl_oai022x1 \REGF/U374  ( .ZN(\REGF/RI_TBAI[9] ), .A(\REGF/n8111 ), .B(
        \REGF/n8225 ), .C(\REGF/n8181 ), .D(\REGF/n8226 ) );
    snl_ao2222x1 \REGF/U542  ( .Z(\REGF/RI_SRDA[15] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[15]), .C(\pgldi[15] ), .D(\REGF/n8210 ), .E(\stream3[15] ), .F(
        \REGF/n8211 ), .G(\pkdptout[15] ), .H(\REGF/n8212 ) );
    snl_and02x1 \REGF/U565  ( .Z(\REGF/RO_LPSAS2156[7] ), .A(
        \REGF/RO_PSASL[9] ), .B(ph_sastlth) );
    snl_invx05 \REGF/U655  ( .ZN(\REGF/n8269 ), .A(ph_stregwt_h) );
    snl_invx05 \REGF/U672  ( .ZN(\REGF/n8193 ), .A(\pgregadrh[7] ) );
    snl_ao01b3x0 \MAIN/U121  ( .Z(\MAIN/*cell*4603/U1/CONTROL1 ), .A(
        \MAIN/n3612 ), .B(wdpr), .C(wspr), .D(ph_lbaovf) );
    snl_ffqrnx1 \MAIN/astregw_tap2_reg  ( .Q(\MAIN/astregw_tap2 ), .D(
        \MAIN/astregw_tap1 ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \LDIS/U148  ( .ZN(\LDIS/n3123 ), .A(\pgld32[23] ) );
    snl_nor02x1 \LDCHK/U34  ( .ZN(LPOUT[3]), .A(\LDCHK/n3231 ), .B(
        \LDCHK/n3235 ) );
    snl_invx05 \LBUS/U688  ( .ZN(\LBUS/n1602 ), .A(\LBUS/n1601 ) );
    snl_muxi21x1 \CODEIF/U299  ( .ZN(\pgfdout[0] ), .A(\CODEIF/n3962 ), .B(
        \CODEIF/n3963 ), .S(mem_cnfg_h) );
    snl_xor2x0 \CODEIF/U309  ( .Z(\CODEIF/n3979 ), .A(CDIN[33]), .B(CDIN[44])
         );
    snl_nand02x1 \ALUIS/U50  ( .ZN(\pgaluinb[2] ), .A(\ALUIS/n3694 ), .B(
        \ALUIS/n3695 ) );
    snl_invx05 \SAEXE/U138  ( .ZN(\SAEXE/n419 ), .A(\SAEXE/n434 ) );
    snl_aoi022x1 \ALUIS/U139  ( .ZN(\ALUIS/n3712 ), .A(\stream4[11] ), .B(
        immbsel), .C(\pk_adb_h[11] ), .D(po_brsel_h) );
    snl_nand02x2 \REGF/U398  ( .ZN(\REGF/n8220 ), .A(ph_sais_h), .B(
        \REGF/n8218 ) );
    snl_ao022x1 \REGF/U419  ( .Z(\REGF/RI_PCOH[14] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[14]), .C(\stream4[46] ), .D(\REGF/n8053 ) );
    snl_oai222x0 \REGF/U442  ( .ZN(\REGF/RI_EACC[23] ), .A(\REGF/n8079 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8080 ), .E(\REGF/n8081 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U459  ( .ZN(\REGF/RI_EACC[6] ), .A(\REGF/n8130 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8131 ), .E(\REGF/n8132 ), 
        .F(\REGF/n8059 ) );
    snl_oai222x0 \REGF/U465  ( .ZN(\REGF/RI_EACC[0] ), .A(\REGF/n8148 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8149 ), .E(\REGF/n8150 ), 
        .F(\REGF/n8059 ) );
    snl_invx05 \REGF/U769  ( .ZN(\REGF/n8170 ), .A(\pgsdprlh[19] ) );
    snl_oai122x0 \CODEIF/U235  ( .ZN(\CODEIF/pfctr415[14] ), .A(\CODEIF/n3864 
        ), .B(\CODEIF/n3908 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3909 ), .E(
        \CODEIF/n3910 ) );
    snl_xnor2x0 \CONS/U244  ( .ZN(\CONS/n520 ), .A(\pk_idcy_h[2] ), .B(
        \pk_indy_h[2] ) );
    snl_xor2x0 \CODEIF/U424  ( .Z(\CODEIF/n3942 ), .A(\CODEIF/n4021 ), .B(
        \CODEIF/n4044 ) );
    snl_invx05 \LBUS/U603  ( .ZN(\LBUS/n1425 ), .A(LDK) );
    snl_ao022x1 \REGF/U817  ( .Z(\REGF/n8244 ), .A(ph_btsrdaselh), .B(
        pk_bitdatah), .C(ph_bdstenh), .D(pk_mpxdh) );
    snl_invx05 \ADOSEL/U49  ( .ZN(\ADOSEL/n4114 ), .A(\pkdptout[8] ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[5]  ( .Q(\CODEIF/pfctr[5] ), .D(
        \CODEIF/pfctr415[5] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_xor2x0 \LDCHK/U98  ( .Z(\LDCHK/n3249 ), .A(\LDCHK/n3310 ), .B(
        \LDCHK/n3295 ) );
    snl_invx05 \LBUS/U624  ( .ZN(\LBUS/n1595 ), .A(\LBUS/EXTSEL ) );
    snl_xnor2x0 \CONS/U174  ( .ZN(\CONS/n653 ), .A(\pgsdprlh[7] ), .B(
        \pk_saco_lh[7] ) );
    snl_nor03x0 \CONS/U153  ( .ZN(\CONS/n726 ), .A(\CONS/n621 ), .B(
        \CONS/n619 ), .C(\CONS/n620 ) );
    snl_invx05 \PDOSEL/U80  ( .ZN(\PDOSEL/n92 ), .A(CDIN[39]) );
    snl_ao222x1 \CODEIF/U209  ( .Z(\CODEIF/n3856 ), .A(PA[18]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[15] ), .E(cif_byte), .F(PDLIN[15]
        ) );
    snl_ao222x1 \CODEIF/U212  ( .Z(\CODEIF/n3859 ), .A(PA[21]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[18] ), .E(cif_byte), .F(PDLIN[18]
        ) );
    snl_xnor2x0 \CODEIF/U382  ( .ZN(\CODEIF/n3951 ), .A(CDIN[43]), .B(CDIN[36]
        ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[16]  ( .Q(\CODEIF/pfctr[16] ), .D(
        \CODEIF/pfctr415[16] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_ao022x1 \REG_2/U132  ( .Z(\ph_cpudout[2] ), .A(\ph_segset_h[2] ), .B(
        seg_cnfg_h), .C(\REG_2/ph_retcnt_h[2] ), .D(ret_cont_h) );
    snl_xnor2x0 \CODEIF/U403  ( .ZN(\CODEIF/n4037 ), .A(CDOUT[56]), .B(CDOUT
        [57]) );
    snl_xnor2x0 \CONS/U263  ( .ZN(\CONS/n744 ), .A(\pk_idcw_h[19] ), .B(
        \pk_indw_h[19] ) );
    snl_xnor2x0 \CODEIF/U399  ( .ZN(\CODEIF/n3993 ), .A(CDIN[1]), .B(CDIN[6])
         );
    snl_xor2x0 \CODEIF/U418  ( .Z(\CODEIF/n3940 ), .A(\CODEIF/n4014 ), .B(
        \CODEIF/n4042 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[3]  ( .Q(CA[3]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3844 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_invx05 \CONS/U278  ( .ZN(\CONS/n551 ), .A(\pgsdprlh[4] ) );
    snl_invx1 \REG_2/U129  ( .ZN(\REG_2/n436 ), .A(\REG_2/n410 ) );
    snl_invx05 \REGF/U755  ( .ZN(\REGF/n8194 ), .A(\pgsdprlh[7] ) );
    snl_invx05 \ADOSEL/U52  ( .ZN(\ADOSEL/n4107 ), .A(\pkdptout[22] ) );
    snl_nor04x0 \LDCHK/U83  ( .ZN(\LDCHK/n3243 ), .A(\pgld32[19] ), .B(
        \pgld32[10] ), .C(\pgld32[20] ), .D(\pgld32[22] ) );
    snl_nor03x0 \CONS/U148  ( .ZN(\CONS/n714 ), .A(\CONS/n612 ), .B(
        \CONS/n610 ), .C(\CONS/n611 ) );
    snl_nand02x1 \PDOSEL/U144  ( .ZN(\PDOSEL/n140 ), .A(CDIN[26]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \REGF/U772  ( .ZN(\REGF/n8176 ), .A(\pgsdprlh[16] ) );
    snl_invx05 \ADOSEL/U75  ( .ZN(\ADOSEL/n4120 ), .A(\pkdptout[10] ) );
    snl_nand02x1 \PDOSEL/U163  ( .ZN(\PDOSEL/n178 ), .A(CDIN[0]), .B(
        \PDOSEL/n119 ) );
    snl_and02x1 \REGF/U830  ( .Z(\REGF/n8219 ), .A(\REGF/n8220 ), .B(
        \REGF/n8221 ) );
    snl_nor02x1 \LBUS/U618  ( .ZN(\LBUS/n1594 ), .A(\LBUS/n1452 ), .B(
        \LBUS/ilt[1] ) );
    snl_oai222x0 \REGF/U480  ( .ZN(\REGF/RI_DPR[13] ), .A(\REGF/n8181 ), .B(
        \REGF/n8160 ), .C(\REGF/n8182 ), .D(\REGF/n8162 ), .E(\REGF/n8111 ), 
        .F(\REGF/n8151 ) );
    snl_ao2222x1 \REGF/U537  ( .Z(\REGF/RI_SRDA[20] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[20]), .C(\pgldi[20] ), .D(\REGF/n8210 ), .E(\stream3[20] ), .F(
        \REGF/n8211 ), .G(\pkdptout[20] ), .H(\REGF/n8212 ) );
    snl_and02x1 \REGF/U559  ( .Z(\REGF/RO_LPSAS2156[1] ), .A(
        \REGF/RO_PSASL[1] ), .B(ph_sastlth) );
    snl_invx05 \REGF/U669  ( .ZN(\REGF/n8123 ), .A(PDLIN[9]) );
    snl_invx05 \CODEIF/U282  ( .ZN(\CODEIF/n3905 ), .A(\CODEIF/pfctr[13] ) );
    snl_xor2x0 \CODEIF/U312  ( .Z(\CODEIF/n3985 ), .A(CDIN[17]), .B(CDIN[16])
         );
    snl_xnor2x0 \LDCHK/U107  ( .ZN(\LDCHK/n3284 ), .A(\pgmuxout[23] ), .B(
        \pgmuxout[21] ) );
    snl_and02x1 \UPIF/U19  ( .Z(\UPIF/n1046 ), .A(WR), .B(\UPIF/ph_accessenh )
         );
    snl_or02x1 \LBUS/U584  ( .Z(ph_piosl_h), .A(\LBUS/PIOSEL_1_Q1249 ), .B(
        ph_ioselh) );
    snl_aoi012x1 \ALUIS/U122  ( .ZN(\ALUIS/n3729 ), .A(\pgldi[19] ), .B(
        srcbsel), .C(allfbsel) );
    snl_muxi21x1 \LDIS/U174  ( .ZN(\LDIS/ldexcl[13] ), .A(\LDIS/n3155 ), .B(
        \LDIS/n3156 ), .S(\LDIS/n3134 ) );
    snl_xor2x0 \CONS/U46  ( .Z(\CONS/n568 ), .A(\pgsdprlh[8] ), .B(
        \pk_saco_lh[8] ) );
    snl_nand02x1 \BLU/U365  ( .ZN(\BLU/n1486 ), .A(\BLU/n1563 ), .B(
        \BLU/n1562 ) );
    snl_invx05 \SAEXE/U123  ( .ZN(\SAEXE/n411 ), .A(\pk_psae_h[5] ) );
    snl_mux21x1 \ALUSHT/U20  ( .Z(\pkdptout[30] ), .A(\ALUSHT/pkshtout[30] ), 
        .B(\ALUSHT/pkaluout[30] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U61  ( .Z(\CONS/n578 ), .A(\pgsdprlh[15] ), .B(
        \CONS/SACO[11] ) );
    snl_and02x2 \UPIF/U7  ( .Z(\ph_pdis_h[6] ), .A(\pk_rread_h[45] ), .B(
        \UPIF/n1046 ) );
    snl_aoi022x1 \LBUS/U693  ( .ZN(\LBUS/n1610 ), .A(\LBUS/n1609 ), .B(
        \pgsadrh[1] ), .C(\LBUS/word32odphase ), .D(\LBUS/n1632 ) );
    snl_ao222x1 \CODEIF/U195  ( .Z(\CODEIF/n3842 ), .A(PA[4]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[1] ), .E(cif_byte), .F(PDLIN[1])
         );
    snl_oai012x1 \PDOSEL/U37  ( .ZN(PDH[53]), .A(\PDOSEL/n107 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_oai022x1 \SAEXE/U104  ( .ZN(ph_wrdsrch), .A(\SAEXE/n413 ), .B(
        \SAEXE/n414 ), .C(\SAEXE/n434 ), .D(\SAEXE/n415 ) );
    snl_invx05 \LDIS/U153  ( .ZN(\LDIS/n3131 ), .A(\pgld32[31] ) );
    snl_oai222x0 \REGF/U607  ( .ZN(\REGF/RI_SPR[22] ), .A(\REGF/n8163 ), .B(
        \REGF/n8220 ), .C(\REGF/n8164 ), .D(\REGF/n8221 ), .E(\REGF/n8084 ), 
        .F(\REGF/n8218 ) );
    snl_xor2x0 \CODEIF/U335  ( .Z(\CODEIF/n4018 ), .A(CDOUT[0]), .B(CDOUT[2])
         );
    snl_xor2x0 \LDCHK/U120  ( .Z(\LDCHK/n3311 ), .A(\LDCHK/n3313 ), .B(
        \LDCHK/n3300 ) );
    snl_nand12x1 \BLU/U342  ( .ZN(\BLU/n1556 ), .A(\poalufnc[4] ), .B(
        \BLU/n1557 ) );
    snl_aoi022x1 \ALUIS/U105  ( .ZN(\ALUIS/n3744 ), .A(\stream4[27] ), .B(
        immbsel), .C(\pk_adb_h[27] ), .D(po_brsel_h) );
    snl_invx05 \REGF/U797  ( .ZN(\REGF/n8074 ), .A(\pkdptout[25] ) );
    snl_nand02x1 \ADOSEL/U90  ( .ZN(\ADOSEL/n4097 ), .A(\pgbluext[2] ), .B(
        \ADOSEL/n4156 ) );
    snl_invx05 \LDCHK/U41  ( .ZN(\LDCHK/n3231 ), .A(ph_ldaoutenhp) );
    snl_nor02x1 \MAIN/U154  ( .ZN(\MAIN/n3629 ), .A(\MAIN/n3623 ), .B(pkaccovf
        ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[2]  ( .Q(\ph_segset_h[2] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[2]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_oai112x0 \PDOSEL/U59  ( .ZN(PDLOUT[14]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n100 ), .C(\PDOSEL/n142 ), .D(\PDOSEL/n143 ) );
    snl_ao022x1 \REGF/U510  ( .Z(\REGF/RI_PCOL[15] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[15]), .C(\stream4[15] ), .D(\REGF/n8209 ) );
    snl_oai222x0 \REGF/U589  ( .ZN(\REGF/RI_ACC[12] ), .A(\REGF/n8112 ), .B(
        \REGF/n8215 ), .C(\REGF/n8113 ), .D(\REGF/n8216 ), .E(\REGF/n8114 ), 
        .F(\REGF/n8217 ) );
    snl_oai222x0 \REGF/U620  ( .ZN(\REGF/RI_SPR[9] ), .A(\REGF/n8189 ), .B(
        \REGF/n8220 ), .C(\REGF/n8190 ), .D(\REGF/n8221 ), .E(\REGF/n8123 ), 
        .F(\REGF/n8218 ) );
    snl_and02x1 \ALUIS/U25  ( .Z(\ALUIS/n3653 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3659 ) );
    snl_xor2x0 \LDCHK/U66  ( .Z(\LDCHK/n3296 ), .A(\pgld32[5] ), .B(
        \LDCHK/pglpinff[0] ) );
    snl_invx05 \CODEIF/U240  ( .ZN(\CODEIF/pgfpcel169 ), .A(\CODEIF/pgfpce_in 
        ) );
    snl_aoi022x1 \ALUIS/U89  ( .ZN(\ALUIS/n3700 ), .A(\stream4[5] ), .B(
        immbsel), .C(\pk_adb_h[5] ), .D(po_brsel_h) );
    snl_invx05 \LBUS/U676  ( .ZN(\LBUS/n1420 ), .A(\LBUS/n1460 ) );
    snl_and08x1 \CONS/U28  ( .Z(ph_iwco_h), .A(\CONS/n338 ), .B(\CONS/n339 ), 
        .C(\CONS/n340 ), .D(\CONS/n341 ), .E(\CONS/n342 ), .F(\CONS/n343 ), 
        .G(\CONS/n344 ), .H(\CONS/n345 ) );
    snl_xor2x0 \CONS/U84  ( .Z(\CONS/n602 ), .A(\pk_idcz_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_xor2x0 \CONS/U101  ( .Z(\CONS/n619 ), .A(\pk_idcx_h[16] ), .B(
        \pk_indx_h[16] ) );
    snl_and02x1 \REG_2/U160  ( .Z(\ph_cpudout[30] ), .A(\ph_segset_h[30] ), 
        .B(seg_cnfg_h) );
    snl_invx05 \CODEIF/U252  ( .ZN(\CODEIF/n3944 ), .A(\CODEIF/wpfcinc ) );
    snl_invx05 \CODEIF/U267  ( .ZN(\CODEIF/n3876 ), .A(PDLIN[3]) );
    snl_xnor2x0 \CONS/U231  ( .ZN(\CONS/n719 ), .A(\pk_idcy_h[10] ), .B(
        \pk_indy_h[10] ) );
    snl_invx05 \BLU/U426  ( .ZN(\BLU/n1546 ), .A(\BLU/n1471 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[12]  ( .Q(\CODEIF/pfctr[12] ), .D(
        \CODEIF/pfctr415[12] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_muxi21x1 \LDIS/U191  ( .ZN(\LDIS/ldexch[19] ), .A(\LDIS/n3146 ), .B(
        \LDIS/n3145 ), .S(\LDIS/n3165 ) );
    snl_and02x1 \CMPX/U9  ( .Z(ph_oprtrs_h), .A(po_oprtrs_h), .B(\CMPX/n1047 )
         );
    snl_nand02x1 \LBUS/U561  ( .ZN(\LBUS/*cell*3982/U148/CONTROL1 ), .A(
        \LBUS/n1400 ), .B(\LBUS/n1401 ) );
    snl_xnor2x0 \CONS/U216  ( .ZN(\CONS/n707 ), .A(\pk_idcz_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_and02x1 \REG_2/U147  ( .Z(\ph_cpudout[17] ), .A(\ph_segset_h[17] ), 
        .B(seg_cnfg_h) );
    snl_nand02x1 \BLU/U380  ( .ZN(\BLU/n1501 ), .A(\BLU/n1568 ), .B(
        \BLU/n1565 ) );
    snl_nand02x1 \BLU/U401  ( .ZN(\BLU/n1510 ), .A(\BLU/n1568 ), .B(
        \BLU/n1563 ) );
    snl_and08x1 \CONS/U126  ( .Z(\CONS/n557 ), .A(\CONS/n657 ), .B(\CONS/n658 
        ), .C(\CONS/n659 ), .D(\CONS/n660 ), .E(\CONS/n661 ), .F(\CONS/n662 ), 
        .G(\CONS/n663 ), .H(\CONS/n656 ) );
    snl_oa012x1 \LBUS/U651  ( .Z(\LBUS/n1433 ), .A(\LBUS/n1423 ), .B(
        \LBUS/n1425 ), .C(\LBUS/n1422 ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[1]  ( .Q(\CODEIF/pfctr[1] ), .D(
        \CODEIF/pfctr415[1] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nand02x1 \LBUS/U664  ( .ZN(\LBUS/n1431 ), .A(\LBUS/n1594 ), .B(
        \LBUS/ilt[5] ) );
    snl_xor2x0 \CONS/U113  ( .Z(\CONS/n631 ), .A(\pk_idcw_h[23] ), .B(
        \pk_indw_h[23] ) );
    snl_xor2x0 \CONS/U96  ( .Z(\CONS/n614 ), .A(\pk_idcy_h[8] ), .B(
        \pk_indy_h[8] ) );
    snl_xnor2x0 \CONS/U223  ( .ZN(\CONS/n711 ), .A(\pk_idcz_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_invx05 \BLU/U434  ( .ZN(\BLU/n1525 ), .A(\BLU/n1519 ) );
    snl_invx05 \CODEIF/U275  ( .ZN(\CODEIF/n3918 ), .A(PDLIN[17]) );
    snl_invx05 \LBUS/U554  ( .ZN(\LBUS/n1393 ), .A(\LBUS/n1392 ) );
    snl_xnor2x0 \CONS/U204  ( .ZN(\CONS/n689 ), .A(\pk_pc_h[6] ), .B(
        \pk_pcs2_h[6] ) );
    snl_and02x1 \REG_2/U155  ( .Z(\ph_cpudout[25] ), .A(\ph_segset_h[25] ), 
        .B(seg_cnfg_h) );
    snl_oa2222x1 \BLU/U413  ( .Z(\BLU/n1516 ), .A(\BLU/n1510 ), .B(\BLU/n1512 
        ), .C(\BLU/n1507 ), .D(\BLU/n1509 ), .E(\BLU/n1504 ), .F(\BLU/n1506 ), 
        .G(\BLU/n1501 ), .H(\BLU/n1503 ) );
    snl_nand13x1 \LBUS/U573  ( .ZN(\LBUS/nlt[1] ), .A(\LBUS/n1427 ), .B(
        \LBUS/n1428 ), .C(\LBUS/n1429 ) );
    snl_invx05 \BLU/U392  ( .ZN(\BLU/n1473 ), .A(\pgld16[13] ) );
    snl_oai222x0 \REGF/U477  ( .ZN(\REGF/RI_DPR[16] ), .A(\REGF/n8175 ), .B(
        \REGF/n8160 ), .C(\REGF/n8176 ), .D(\REGF/n8162 ), .E(\REGF/n8102 ), 
        .F(\REGF/n8151 ) );
    snl_oai222x0 \REGF/U492  ( .ZN(\REGF/RI_DPR[1] ), .A(\REGF/n8205 ), .B(
        \REGF/n8160 ), .C(\REGF/n8206 ), .D(\REGF/n8162 ), .E(\REGF/n8147 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U502  ( .Z(\REGF/RI_PCOL[23] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[23]), .C(\stream4[23] ), .D(\REGF/n8209 ) );
    snl_ao022x1 \REGF/U525  ( .Z(\REGF/RI_PCOL[0] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[0]), .C(\stream4[0] ), .D(\REGF/n8209 ) );
    snl_oai222x0 \REGF/U615  ( .ZN(\REGF/RI_SPR[14] ), .A(\REGF/n8179 ), .B(
        \REGF/n8220 ), .C(\REGF/n8180 ), .D(\REGF/n8221 ), .E(\REGF/n8108 ), 
        .F(\REGF/n8218 ) );
    snl_invx05 \REGF/U729  ( .ZN(\REGF/n8067 ), .A(\pgldi[27] ) );
    snl_muxi21x1 \LDIS/U183  ( .ZN(\LDIS/ldexch[27] ), .A(\LDIS/n3160 ), .B(
        \LDIS/n3159 ), .S(\LDIS/n3165 ) );
    snl_sffqqnx1 \LBUS/pdchken_reg  ( .QN(\LBUS/n1391 ), .D(\LBUS/temp[3] ), 
        .SD(1'b0), .SE(ph_lbwrh), .CP(SCLK) );
    snl_and08x1 \CONS/U134  ( .Z(\CONS/n646 ), .A(\CONS/n675 ), .B(\CONS/n676 
        ), .C(\CONS/n677 ), .D(\CONS/n678 ), .E(\CONS/n679 ), .F(\CONS/n680 ), 
        .G(\CONS/n681 ), .H(\CONS/n674 ) );
    snl_nand02x1 \PDOSEL/U138  ( .ZN(\PDOSEL/n156 ), .A(CDIN[6]), .B(
        \PDOSEL/n119 ) );
    snl_invx05 \REGF/U785  ( .ZN(\REGF/n8128 ), .A(\pkdptout[7] ) );
    snl_muxi21x1 \LDCHK/U53  ( .ZN(\LDCHK/lpex[2] ), .A(\LDCHK/n3275 ), .B(
        \LDCHK/n3276 ), .S(\LDCHK/n3274 ) );
    snl_oai012x1 \LBUS/U643  ( .ZN(\LBUS/n1399 ), .A(\LBUS/n1451 ), .B(
        \LBUS/n1463 ), .C(\LBUS/n1398 ) );
    snl_ffqrnx1 \SAEXE/ph_lmterr_h_reg  ( .Q(phlmterr_h), .D(
        \SAEXE/*cell*3651/U4/CONTROL1 ), .RN(n10735), .CP(SCLK) );
    snl_nand02x1 \ADOSEL/U82  ( .ZN(\ADOSEL/n4115 ), .A(\pgbluext[8] ), .B(
        \ADOSEL/n4156 ) );
    snl_aoi022x1 \MAIN/U146  ( .ZN(\MAIN/n3630 ), .A(\MAIN/ph_rdwr1selh ), .B(
        wonly1), .C(\MAIN/ph_rdwr2selh ), .D(wonly2) );
    snl_xnor2x0 \CONS/U198  ( .ZN(\CONS/n679 ), .A(\pk_pc_h[4] ), .B(
        \pk_pcs2_h[4] ) );
    snl_nand02x1 \CODEIF/U349  ( .ZN(\CODEIF/n3919 ), .A(\CODEIF/pgctrinc[17] 
        ), .B(\CODEIF/n3945 ) );
    snl_and02x1 \ALUIS/U10  ( .Z(\ALUIS/n3643 ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3660 ) );
    snl_ao02b2x1 \REGF/U632  ( .Z(\REGF/RI_STAT[3] ), .A(\REGF/n8223 ), .B(
        \REGF/n8096 ), .C(\REGF/n8224 ), .D(oltff) );
    snl_nand02x1 \ALUIS/U37  ( .ZN(\pgaluina[21] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3679 ) );
    snl_aoi0b12x0 \BLU/U319  ( .ZN(\BLU/n1519 ), .A(\pk_stat_h[0] ), .B(
        accasel), .C(\BLU/n1520 ) );
    snl_invx05 \CODEIF/U290  ( .ZN(\CODEIF/n3865 ), .A(\CODEIF/pfctr[0] ) );
    snl_invx05 \MAIN/U161  ( .ZN(ph_ciwt_h), .A(\MAIN/n3614 ) );
    snl_xor2x0 \LDCHK/U74  ( .Z(\LDCHK/n3264 ), .A(\LDCHK/n3301 ), .B(
        \LDCHK/n3302 ) );
    snl_xnor2x0 \LDCHK/U115  ( .ZN(\LDCHK/n3292 ), .A(\pgmuxout[4] ), .B(
        \pgmuxout[2] ) );
    snl_ao022x1 \LDIS/U108  ( .Z(\pgldi[5] ), .A(ph_word32_h), .B(\pgld32[5] ), 
        .C(\pgld16[5] ), .D(ph_word16_h) );
    snl_invx05 \CMPX/U19  ( .ZN(\CMPX/n1050 ), .A(phadrdech) );
    snl_nor02x1 \LBUS/U596  ( .ZN(\LBUS/n1447 ), .A(ph_word32_h), .B(
        ph_word16_h) );
    snl_sffqenrnx1 \REG_2/RETCNT_reg[7]  ( .Q(\REG_2/RETCNT[7] ), .D(
        \REG_2/ph_retcnt_h[7] ), .EN(\REG_2/n517 ), .RN(\REG_2/n435 ), .SD(
        \REG_2/ncnt3[1] ), .SE(ph_d76lth), .CP(SCLK) );
    snl_xor2x0 \CODEIF/U300  ( .Z(\CODEIF/n3947 ), .A(\CODEIF/n3964 ), .B(
        \CODEIF/n3965 ) );
    snl_nand02x1 \BLU/U377  ( .ZN(\BLU/n1498 ), .A(\BLU/n1569 ), .B(
        \BLU/n1563 ) );
    snl_xor2x0 \CODEIF/U327  ( .Z(\CODEIF/n4006 ), .A(CDOUT[41]), .B(CDOUT[32]
        ) );
    snl_nand02x1 \ALUIS/U59  ( .ZN(\pgaluinb[11] ), .A(\ALUIS/n3712 ), .B(
        \ALUIS/n3713 ) );
    snl_aoi012x1 \ALUIS/U130  ( .ZN(\ALUIS/n3721 ), .A(\pgldi[15] ), .B(
        srcbsel), .C(allfbsel) );
    snl_or02x1 \MAIN/U128  ( .Z(\MAIN/astregw_inhibith ), .A(
        \MAIN/astregw_tap2 ), .B(\MAIN/astregw_tap1 ) );
    snl_oai012x1 \LDIS/U141  ( .ZN(\pgldi[27] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3127 ), .C(\LDIS/n3115 ) );
    snl_muxi21x1 \LDIS/U166  ( .ZN(\LDIS/ldexcl[6] ), .A(\LDIS/n3139 ), .B(
        \LDIS/n3140 ), .S(\LDIS/n3134 ) );
    snl_mux21x1 \ALUSHT/U15  ( .Z(\pkdptout[6] ), .A(\ALUSHT/pkshtout[6] ), 
        .B(\ALUSHT/pkaluout[6] ), .S(\ALUSHT/n3112 ) );
    snl_xor2x0 \CONS/U54  ( .Z(\CONS/n564 ), .A(\pgsdprlh[12] ), .B(
        \CONS/SACO[8] ) );
    snl_nand13x1 \SAEXE/U131  ( .ZN(\SAEXE/n414 ), .A(\pk_psae_h[1] ), .B(
        \SAEXE/n429 ), .C(\pk_psae_h[0] ) );
    snl_mux21x1 \ALUSHT/U32  ( .Z(\pkdptout[1] ), .A(\ALUSHT/pkshtout[1] ), 
        .B(\ALUSHT/pkaluout[1] ), .S(\ALUSHT/n3112 ) );
    snl_and34x0 \SAEXE/U116  ( .Z(phadrdech), .A(\pk_psae_h[7] ), .B(
        \pk_psae_h[2] ), .C(\SAEXE/n413 ), .D(\pk_psae_h[3] ) );
    snl_and02x1 \LBUS/U681  ( .Z(\LBUS/n1411 ), .A(\LBUS/n1610 ), .B(
        \LBUS/n1608 ) );
    snl_xor2x0 \CONS/U73  ( .Z(\CONS/n591 ), .A(\pk_pc_h[5] ), .B(
        \pk_pcs1_h[5] ) );
    snl_oai012x1 \PDOSEL/U25  ( .ZN(PDH[41]), .A(\PDOSEL/n95 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[12]  ( .Q(CA[12]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3853 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_aoi022x1 \ALUIS/U117  ( .ZN(\ALUIS/n3732 ), .A(\stream4[21] ), .B(
        immbsel), .C(\pk_adb_h[21] ), .D(po_brsel_h) );
    snl_nor02x1 \BLU/U350  ( .ZN(\BLU/n1565 ), .A(\BLU/n1564 ), .B(\BLU/n1560 
        ) );
    snl_invx05 \REGF/U805  ( .ZN(\REGF/n8095 ), .A(\pkdptout[18] ) );
    snl_oai122x0 \ADOSEL/U40  ( .ZN(\pgmuxout[29] ), .A(\ADOSEL/n4137 ), .B(
        \ADOSEL/n4129 ), .C(\ADOSEL/n4138 ), .D(\ADOSEL/n4128 ), .E(
        \ADOSEL/n4152 ) );
    snl_invx05 \PDOSEL/U89  ( .ZN(\PDOSEL/n110 ), .A(CDIN[56]) );
    snl_nand02x1 \PDOSEL/U156  ( .ZN(\PDOSEL/n150 ), .A(CDIN[16]), .B(
        \PDOSEL/n119 ) );
    snl_oai222x0 \REGF/U450  ( .ZN(\REGF/RI_EACC[15] ), .A(\REGF/n8103 ), .B(
        \REGF/n8055 ), .C(\REGF/n8056 ), .D(\REGF/n8104 ), .E(\REGF/n8105 ), 
        .F(\REGF/n8059 ) );
    snl_invx05 \REGF/U747  ( .ZN(\REGF/n8106 ), .A(\pgldi[14] ) );
    snl_invx05 \REGF/U760  ( .ZN(\REGF/n8201 ), .A(\pgregadrh[3] ) );
    snl_invx05 \ADOSEL/U67  ( .ZN(\ADOSEL/n4095 ), .A(\pkdptout[18] ) );
    snl_invx05 \LDCHK/U91  ( .ZN(\LDCHK/n3276 ), .A(LPIN[0]) );
    snl_mux21x2 \SHTCD/U11  ( .Z(\phshtd[3] ), .A(\pgld16[3] ), .B(
        \stream4[3] ), .S(immbsel) );
    snl_nand04x0 \REGF/U822  ( .ZN(\REGF/n8235 ), .A(pk_sign_h), .B(
        \REGF/RO_ACC[30] ), .C(\REGF/RO_ACC[25] ), .D(\REGF/RO_ACC[26] ) );
    snl_oai2222x0 \REGF/U366  ( .ZN(\REGF/RI_SRA12M[3] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8141 ), .C(\REGF/n8139 ), .D(\REGF/n8051 ), .E(\REGF/n8229 ), 
        .F(\REGF/n8201 ), .G(\REGF/n8230 ), .H(\REGF/n8202 ) );
    snl_ao2222x1 \REGF/U550  ( .Z(\REGF/RI_SRDA[7] ), .A(\ph_pdis_h[9] ), .B(
        PDLIN[7]), .C(\pgldi[7] ), .D(\REGF/n8210 ), .E(\stream3[7] ), .F(
        \REGF/n8211 ), .G(\pkdptout[7] ), .H(\REGF/n8212 ) );
    snl_nand02x1 \ADOSEL/U103  ( .ZN(\ADOSEL/n4141 ), .A(\pgbluext[2] ), .B(
        \ADOSEL/n4156 ) );
    snl_ao222x1 \CODEIF/U200  ( .Z(\CODEIF/n3847 ), .A(PA[9]), .B(cif_cont), 
        .C(\CODEIF/n3929 ), .D(\CODEIF/pfctr[6] ), .E(cif_byte), .F(PDLIN[6])
         );
    snl_oai122x0 \CODEIF/U227  ( .ZN(\CODEIF/pfctr415[6] ), .A(\CODEIF/n3864 ), 
        .B(\CODEIF/n3884 ), .C(\CODEIF/n3867 ), .D(\CODEIF/n3885 ), .E(
        \CODEIF/n3886 ) );
    snl_sffqenrnx1 \LDCHK/pglpinff_reg[1]  ( .Q(\LDCHK/pglpinff[1] ), .D(1'b0), 
        .EN(1'b1), .RN(n10733), .SD(\LDCHK/lpex[1] ), .SE(ph_lpdilth), .CP(
        SCLK) );
    snl_nand03x0 \LBUS/U611  ( .ZN(\LBUS/n1461 ), .A(\LBUS/ilt[1] ), .B(LASOUT
        ), .C(\LBUS/n1460 ) );
    snl_xnor2x0 \CONS/U256  ( .ZN(\CONS/n733 ), .A(\pk_idcx_h[11] ), .B(
        \pk_indx_h[11] ) );
    snl_invx05 \BLU/U441  ( .ZN(pk_mpxdh), .A(\BLU/n1464 ) );
    snl_oai222x0 \CONS/U166  ( .ZN(\CONS/n640 ), .A(\CONS/n545 ), .B(
        \CONS/n549 ), .C(\CONS/n539 ), .D(\CONS/n547 ), .E(\CONS/n550 ), .F(
        \CONS/n559 ) );
    snl_nor03x0 \LBUS/U636  ( .ZN(\LBUS/n1601 ), .A(ph_errtendh), .B(
        \LBUS/MMBSEL ), .C(\LBUS/OBMSEL ) );
    snl_nor04x0 \CONS/U141  ( .ZN(\CONS/n643 ), .A(\CONS/n699 ), .B(
        \CONS/n596 ), .C(\CONS/n594 ), .D(\CONS/n595 ) );
    snl_invx05 \PDOSEL/U92  ( .ZN(\PDOSEL/n107 ), .A(CDIN[53]) );
    snl_xor2x0 \CODEIF/U390  ( .Z(\CODEIF/n4033 ), .A(\CODEIF/n3982 ), .B(
        \CODEIF/n3986 ) );
    snl_xnor2x0 \CONS/U271  ( .ZN(\CONS/n745 ), .A(\pk_idcw_h[17] ), .B(
        \pk_indw_h[17] ) );
    snl_xor2x0 \CODEIF/U411  ( .Z(\CODEIF/n4040 ), .A(\CODEIF/n4005 ), .B(
        \CODEIF/n4001 ) );
    snl_nand02x1 \ALUIS/U65  ( .ZN(\pgaluinb[17] ), .A(\ALUIS/n3724 ), .B(
        \ALUIS/n3725 ) );
    snl_oai022x1 \REGF/U647  ( .ZN(\REGF/RI_TBAI[7] ), .A(\REGF/n8225 ), .B(
        \REGF/n8117 ), .C(\REGF/n8226 ), .D(\REGF/n8185 ) );
    snl_invx05 \REGF/U660  ( .ZN(\REGF/n8181 ), .A(\pgregadrh[13] ) );
    snl_oai122x0 \MAIN/U133  ( .ZN(\MAIN/reg_enable ), .A(saenabl1), .B(
        \MAIN/n3627 ), .C(saenabl2), .D(\MAIN/n3628 ), .E(\MAIN/n3629 ) );
    snl_mux21x1 \ALUSHT/U29  ( .Z(\pkdptout[22] ), .A(\ALUSHT/pkshtout[22] ), 
        .B(\ALUSHT/pkaluout[22] ), .S(\ALUSHT/n3112 ) );
    snl_sffqenrnx1 \LBUS/ph_selldl_reg  ( .Q(ph_selldl), .D(1'b0), .EN(1'b1), 
        .RN(n10734), .SD(\LBUS/n1632 ), .SE(\LBUS/*cell*3982/U188/CONTROL1 ), 
        .CP(SCLK) );
    snl_xor2x0 \CONS/U68  ( .Z(\CONS/n586 ), .A(\pk_pc_h[2] ), .B(
        \pk_pcs2_h[2] ) );
    snl_oai012x1 \PDOSEL/U19  ( .ZN(PDH[35]), .A(\PDOSEL/n79 ), .B(
        \PDOSEL/n75 ), .C(\PDOSEL/n76 ) );
    snl_nand02x1 \ALUIS/U42  ( .ZN(\pgaluina[26] ), .A(\ALUIS/n3657 ), .B(
        \ALUIS/n3684 ) );
    snl_and02x1 \UPIF/U10  ( .Z(\ph_pdis_h[10] ), .A(\pk_rread_h[38] ), .B(
        \UPIF/n1046 ) );
    snl_oai2222x0 \REGF/U383  ( .ZN(\REGF/RI_SRA12M[11] ), .A(\REGF/n8228 ), 
        .B(\REGF/n8117 ), .C(\REGF/n8115 ), .D(\REGF/n8051 ), .E(\REGF/n8185 ), 
        .F(\REGF/n8229 ), .G(\REGF/n8230 ), .H(\REGF/n8186 ) );
    snl_nand02x2 \REGF/U402  ( .ZN(\REGF/n8162 ), .A(po_ptrsel_h), .B(
        \REGF/n8151 ) );
    snl_oai222x0 \REGF/U489  ( .ZN(\REGF/RI_DPR[4] ), .A(\REGF/n8199 ), .B(
        \REGF/n8160 ), .C(\REGF/n8200 ), .D(\REGF/n8162 ), .E(\REGF/n8138 ), 
        .F(\REGF/n8151 ) );
    snl_ao022x1 \REGF/U519  ( .Z(\REGF/RI_PCOL[6] ), .A(\ph_pdis_h[6] ), .B(
        PDLIN[6]), .C(\stream4[6] ), .D(\REGF/n8209 ) );
    snl_oai222x0 \REGF/U577  ( .ZN(\REGF/RI_ACC[24] ), .A(\REGF/n8076 ), .B(
        \REGF/n8215 ), .C(\REGF/n8077 ), .D(\REGF/n8216 ), .E(\REGF/n8078 ), 
        .F(\REGF/n8217 ) );
    snl_sffqenrnx1 \REG_2/ph_segset_h_reg[6]  ( .Q(\ph_segset_h[6] ), .D(1'b0), 
        .EN(1'b1), .RN(\REG_2/n436 ), .SD(PDLIN[6]), .SE(seg_config_wr), .CP(
        SCLK) );
    snl_oai222x0 \REGF/U629  ( .ZN(\REGF/RI_SPR[0] ), .A(\REGF/n8207 ), .B(
        \REGF/n8220 ), .C(\REGF/n8208 ), .D(\REGF/n8221 ), .E(\REGF/n8150 ), 
        .F(\REGF/n8218 ) );
    snl_ao022x1 \LDIS/U113  ( .Z(\pgld16[7] ), .A(ph_selldl), .B(\pgld32[7] ), 
        .C(ph_selldh), .D(\pgld32[23] ) );
    snl_and02x1 \PDOSEL/U77  ( .Z(\PDOSEL/n119 ), .A(\PDOSEL/n224 ), .B(
        code_area_h) );
    snl_xnor2x0 \CODEIF/U375  ( .ZN(\CODEIF/n3948 ), .A(CDIN[51]), .B(CDIN[59]
        ) );
    snl_nand02x1 \ALUIS/U145  ( .ZN(\ALUIS/n3666 ), .A(\pk_ada_h[8] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U223  ( .ZN(\LDIS/n3153 ), .A(LIN[14]) );
    snl_oai022x1 \BLU/U302  ( .ZN(\pkbludgh[14] ), .A(\BLU/n1464 ), .B(
        \BLU/n1468 ), .C(\BLU/n1469 ), .D(\BLU/n1470 ) );
    snl_oai222x0 \REGF/U592  ( .ZN(\REGF/RI_ACC[9] ), .A(\REGF/n8121 ), .B(
        \REGF/n8215 ), .C(\REGF/n8122 ), .D(\REGF/n8216 ), .E(\REGF/n8123 ), 
        .F(\REGF/n8217 ) );
    snl_invx05 \REGF/U732  ( .ZN(\REGF/n8072 ), .A(PDLIN[26]) );
    snl_nand02x1 \ADOSEL/U99  ( .ZN(\ADOSEL/n4144 ), .A(\pgbluext[5] ), .B(
        \ADOSEL/n4156 ) );
    snl_nand02x1 \CODEIF/U352  ( .ZN(\CODEIF/n3910 ), .A(\CODEIF/pgctrinc[14] 
        ), .B(\CODEIF/n3945 ) );
    snl_nor02x1 \BLU/U325  ( .ZN(\BLU/n1493 ), .A(\BLU/n1535 ), .B(\BLU/n1536 
        ) );
    snl_ffqrnx1 \CODEIF/pfctr_reg[8]  ( .Q(\CODEIF/pfctr[8] ), .D(
        \CODEIF/pfctr415[8] ), .RN(\CODEIF/n3861 ), .CP(SCLK) );
    snl_nand02x1 \ALUIS/U162  ( .ZN(\ALUIS/n3679 ), .A(\pk_ada_h[21] ), .B(
        po_arsel_h) );
    snl_invx05 \LDIS/U204  ( .ZN(\LDIS/n3144 ), .A(LIN[20]) );
    snl_ao022x1 \CMPX/U25  ( .Z(ph_lmterr_h), .A(phlmterr_h), .B(ph_saexe_sth), 
        .C(phlmterrh), .D(\CMPX/n1047 ) );
    snl_xor2x0 \LDCHK/U48  ( .Z(\LDCHK/n3254 ), .A(\LDCHK/n3264 ), .B(
        \LDCHK/n3265 ) );
    snl_oai012x1 \LDIS/U134  ( .ZN(\pgldi[20] ), .A(\LDIS/n3113 ), .B(
        \LDIS/n3120 ), .C(\LDIS/n3115 ) );
    snl_xnor2x0 \CONS/U183  ( .ZN(\CONS/n661 ), .A(\pgsdprlh[12] ), .B(
        \pk_saco_lh[12] ) );
    snl_oai112x0 \PDOSEL/U50  ( .ZN(PDLOUT[11]), .A(\PDOSEL/n114 ), .B(
        \PDOSEL/n97 ), .C(\PDOSEL/n126 ), .D(\PDOSEL/n127 ) );
    snl_invx05 \LBUS/U658  ( .ZN(\LBUS/*cell*3982/U31/CONTROL1 ), .A(
        \LBUS/n1413 ) );
    snl_oai122x0 \ADOSEL/U35  ( .ZN(\pgmuxout[24] ), .A(\ADOSEL/n4114 ), .B(
        \ADOSEL/n4137 ), .C(\ADOSEL/n4113 ), .D(\ADOSEL/n4138 ), .E(
        \ADOSEL/n4147 ) );
    snl_invx05 \LDIS/U198  ( .ZN(\LDIS/n3150 ), .A(LIN[17]) );
    snl_aoi112x0 \PDOSEL/U123  ( .ZN(\PDOSEL/n121 ), .A(\pgfdout[1] ), .B(
        \PDOSEL/n226 ), .C(\ph_cpudout[1] ), .D(\pk_pdo_h[1] ) );
    snl_ao022x1 \REGF/U425  ( .Z(\REGF/RI_PCOH[8] ), .A(\ph_pdis_h[5] ), .B(
        PDLIN[8]), .C(\stream4[40] ), .D(\REGF/n8053 ) );
    snl_nand02x1 \LBUS/U568  ( .ZN(\LBUS/*cell*3982/U185/CONTROL1 ), .A(
        \LBUS/n1405 ), .B(\LBUS/n1413 ) );
    snl_nand13x1 \BLU/U389  ( .ZN(\BLU/n1547 ), .A(\BLU/n1545 ), .B(
        \BLU/n1465 ), .C(\BLU/n1474 ) );
    snl_muxi21x1 \BLU/U408  ( .ZN(oebacc), .A(\BLU/n1580 ), .B(\BLU/n1581 ), 
        .S(ph_shelter_h) );
    snl_invx05 \REGF/U685  ( .ZN(\REGF/n8135 ), .A(PDLIN[5]) );
    snl_and12x1 \REGF/U715  ( .Z(\REGF/n8210 ), .A(\ph_pdis_h[9] ), .B(
        ph_wdsrdaselh) );
    snl_invx05 \CODEIF/U249  ( .ZN(\CODEIF/n3927 ), .A(\CODEIF/write_prtect )
         );
    snl_sffqenrnx1 \CODEIF/pgfadrh_reg[7]  ( .Q(CA[7]), .D(1'b0), .EN(1'b1), 
        .RN(\CODEIF/n3862 ), .SD(\CODEIF/n3848 ), .SE(\CODEIF/fadren ), .CP(
        SCLK) );
    snl_aoi012x1 \ALUIS/U80  ( .ZN(\ALUIS/n3709 ), .A(srcbsel), .B(\pgldi[9] ), 
        .C(allfbsel) );
    snl_xnor2x0 \CONS/U238  ( .ZN(\CONS/n723 ), .A(\pk_idcy_h[21] ), .B(
        \pk_indy_h[21] ) );
    snl_oai122x0 \ADOSEL/U12  ( .ZN(\pgmuxout[1] ), .A(\ADOSEL/n4087 ), .B(
        \ADOSEL/n4092 ), .C(\ADOSEL/n4089 ), .D(\ADOSEL/n4093 ), .E(
        \ADOSEL/n4094 ) );
    snl_xor2x0 \CONS/U108  ( .Z(\CONS/n626 ), .A(\pk_idcx_h[18] ), .B(
        \pk_indx_h[18] ) );
    snl_invx05 \PDOSEL/U104  ( .ZN(\PDOSEL/n96 ), .A(CDIN[42]) );
    snl_and34x1 \MCD/insdec_1/U163  ( .Z(po_ldis_h), .A(\MCD/insdec_1/n4196 ), 
        .B(\MCD/insdec_1/n4197 ), .C(\MCD/insdec_1/n4169 ), .D(
        \MCD/insdec_1/n4195 ) );
    snl_aoi013x2 \MCD/insdec_1/U165  ( .ZN(\MCD/insdec_1/n4184 ), .A(
        \MCD/insdec_1/n4223 ), .B(\MCD/insdec_1/n4182 ), .C(
        \MCD/insdec_1/n4241 ), .D(\MCD/insdec_1/n4213 ) );
    snl_nor04x8 \MCD/insdec_1/U166  ( .ZN(immbsel), .A(ph_saexe_sth), .B(
        \stream4[47] ), .C(\MCD/insdec_1/n4184 ), .D(\MCD/insdec_1/n4185 ) );
    snl_oai112x0 \MCD/insdec_1/U198  ( .ZN(\MCD/insdec_1/n4202 ), .A(
        \MCD/insdec_1/n4217 ), .B(\MCD/insdec_1/n4218 ), .C(
        \MCD/insdec_1/n4219 ), .D(\MCD/insdec_1/n4220 ) );
    snl_nor02x1 \MCD/insdec_1/U204  ( .ZN(\MCD/insdec_1/n4230 ), .A(
        \MCD/insdec_1/n4203 ), .B(\MCD/insdec_1/n4231 ) );
    snl_nor02x1 \MCD/insdec_1/U223  ( .ZN(\MCD/insdec_1/n4229 ), .A(
        pk_pcon31_h), .B(\MCD/insdec_1/n4250 ) );
    snl_oai233x1 \MCD/insdec_1/U167  ( .ZN(\poalufnc[4] ), .A(
        \MCD/insdec_1/n4158 ), .B(\MCD/insdec_1/n4159 ), .C(
        \MCD/insdec_1/n4160 ), .D(\MCD/insdec_1/n4161 ), .E(\stream4[38] ), 
        .F(\stream4[37] ), .G(\MCD/insdec_1/n4162 ), .H(\MCD/insdec_1/n4163 )
         );
    snl_ao022x2 \MCD/insdec_1/U168  ( .Z(srcbsel), .A(ph_srcsl_h), .B(
        ph_saexe_sth), .C(\MCD/insdec_1/n4195 ), .D(\MCD/insdec_1/n4165 ) );
    snl_nor03x4 \MCD/insdec_1/U174  ( .ZN(accbsel), .A(\MCD/insdec_1/n4184 ), 
        .B(ph_saexe_sth), .C(\MCD/insdec_1/n4237 ) );
    snl_nor03x0 \MCD/insdec_1/U183  ( .ZN(ebaccsel), .A(\MCD/insdec_1/n4178 ), 
        .B(\MCD/insdec_1/n4179 ), .C(\MCD/insdec_1/n4180 ) );
    snl_and03x1 \MCD/insdec_1/U256  ( .Z(\MCD/insdec_1/n4268 ), .A(
        \MCD/insdec_1/n4229 ), .B(\MCD/insdec_1/n4254 ), .C(
        \MCD/insdec_1/n4239 ) );
    snl_nand02x1 \MCD/insdec_1/U271  ( .ZN(\MCD/insdec_1/n4219 ), .A(
        \MCD/insdec_1/n4278 ), .B(\MCD/insdec_1/n4253 ) );
    snl_invx05 \MCD/insdec_1/U294  ( .ZN(\MCD/insdec_1/n4206 ), .A(
        \MCD/insdec_1/n4161 ) );
    snl_and02x1 \MCD/insdec_1/U304  ( .Z(\MCD/insdec_1/n4167 ), .A(
        \stream4[38] ), .B(\MCD/insdec_1/n4163 ) );
    snl_aoi022x1 \MCD/insdec_1/U191  ( .ZN(\MCD/insdec_1/n4200 ), .A(
        ph_piosl_h), .B(\pk_stat_h[18] ), .C(\MCD/insdec_1/bacc ), .D(
        \MCD/insdec_1/ciff ) );
    snl_invx05 \MCD/insdec_1/U238  ( .ZN(\MCD/insdec_1/n4163 ), .A(
        \stream4[39] ) );
    snl_nand02x1 \MCD/insdec_1/U286  ( .ZN(\MCD/insdec_1/n4186 ), .A(
        \MCD/insdec_1/n4192 ), .B(\MCD/insdec_1/n4165 ) );
    snl_aoi022x1 \MCD/insdec_1/U316  ( .ZN(\MCD/insdec_1/n4257 ), .A(
        \MCD/insdec_1/n4268 ), .B(\stream4[33] ), .C(\MCD/insdec_1/n4269 ), 
        .D(\MCD/insdec_1/n4247 ) );
    snl_ffqrnx1 \MCD/insdec_1/ciff_reg  ( .Q(\MCD/insdec_1/ciff ), .D(pk_ciffh
        ), .RN(n10733), .CP(SCLK) );
    snl_nor02x1 \MCD/insdec_1/U211  ( .ZN(\MCD/insdec_1/n4223 ), .A(
        \stream4[59] ), .B(\stream4[58] ) );
    snl_invx05 \MCD/insdec_1/U216  ( .ZN(\MCD/insdec_1/n4180 ), .A(
        \stream4[40] ) );
    snl_oai112x0 \MCD/insdec_1/U231  ( .ZN(\MCD/insdec_1/n4224 ), .A(
        \MCD/insdec_1/n4252 ), .B(\MCD/insdec_1/n4217 ), .C(
        \MCD/insdec_1/n4215 ), .D(\MCD/insdec_1/n4216 ) );
    snl_nor02x1 \MCD/insdec_1/U244  ( .ZN(\MCD/insdec_1/n4222 ), .A(
        \stream4[50] ), .B(\stream4[51] ) );
    snl_nor02x1 \MCD/insdec_1/U263  ( .ZN(\MCD/insdec_1/n4242 ), .A(
        \stream4[41] ), .B(\MCD/insdec_1/n4180 ) );
    snl_invx05 \MCD/insdec_1/U278  ( .ZN(\MCD/insdec_1/n4159 ), .A(
        \MCD/insdec_1/n4214 ) );
    snl_nand02x1 \MCD/insdec_1/U236  ( .ZN(\MCD/insdec_1/n4158 ), .A(
        \MCD/insdec_1/n4170 ), .B(\MCD/insdec_1/n4262 ) );
    snl_ao112x2 \MCD/insdec_1/U169  ( .Z(po_brsel_h), .A(ph_dregsl_h), .B(
        ph_saexe_sth), .C(eaccbsel), .D(accbsel) );
    snl_nor03x2 \MCD/insdec_1/U172  ( .ZN(exetype1), .A(\stream4[56] ), .B(
        \stream4[59] ), .C(\MCD/insdec_1/n4245 ) );
    snl_nor03x4 \MCD/insdec_1/U173  ( .ZN(allfbsel), .A(\MCD/insdec_1/n4181 ), 
        .B(ph_saexe_sth), .C(\MCD/insdec_1/n4182 ) );
    snl_invx05 \MCD/insdec_1/U243  ( .ZN(\MCD/insdec_1/n4165 ), .A(
        ph_saexe_sth) );
    snl_nand02x1 \MCD/insdec_1/U258  ( .ZN(\MCD/insdec_1/n4270 ), .A(
        \MCD/insdec_1/ciff ), .B(\stream4[32] ) );
    snl_nor02x1 \MCD/insdec_1/U264  ( .ZN(\MCD/insdec_1/n4243 ), .A(
        \stream4[43] ), .B(\MCD/insdec_1/n4265 ) );
    snl_nor02x1 \MCD/insdec_1/U184  ( .ZN(allfasel), .A(ph_saexe_sth), .B(
        \MCD/insdec_1/n4183 ) );
    snl_aoi012x1 \MCD/insdec_1/U196  ( .ZN(\MCD/insdec_1/n4209 ), .A(
        \MCD/insdec_1/n4210 ), .B(\MCD/insdec_1/n4211 ), .C(
        \MCD/insdec_1/n4212 ) );
    snl_and23x0 \MCD/insdec_1/U281  ( .Z(srctype1), .A(\stream4[53] ), .B(
        \stream4[54] ), .C(\stream4[52] ) );
    snl_invx05 \MCD/insdec_1/U311  ( .ZN(\MCD/insdec_1/n4274 ), .A(
        \MCD/insdec_1/n4276 ) );
    snl_nand03x0 \MCD/insdec_1/U197  ( .ZN(\MCD/insdec_1/n4213 ), .A(
        \MCD/insdec_1/n4214 ), .B(\MCD/insdec_1/n4215 ), .C(
        \MCD/insdec_1/n4216 ) );
    snl_nor02x1 \MCD/insdec_1/U203  ( .ZN(\MCD/insdec_1/n4228 ), .A(
        \stream4[32] ), .B(\MCD/insdec_1/n4229 ) );
    snl_invx05 \MCD/insdec_1/U218  ( .ZN(\MCD/insdec_1/n4247 ), .A(
        \stream4[33] ) );
    snl_invx05 \MCD/insdec_1/U293  ( .ZN(\MCD/insdec_1/n4264 ), .A(
        \MCD/insdec_1/n4222 ) );
    snl_invx05 \MCD/insdec_1/U303  ( .ZN(\MCD/insdec_1/n4173 ), .A(
        \poalufnc[3] ) );
    snl_nand03x0 \MCD/insdec_1/U251  ( .ZN(\MCD/insdec_1/n4178 ), .A(
        \MCD/insdec_1/n4245 ), .B(\MCD/insdec_1/n4165 ), .C(
        \MCD/insdec_1/n4199 ) );
    snl_nand02x1 \MCD/insdec_1/U276  ( .ZN(\MCD/insdec_1/n4215 ), .A(
        \MCD/insdec_1/n4253 ), .B(stage_b) );
    snl_nand02x1 \MCD/insdec_1/U224  ( .ZN(\MCD/insdec_1/n4251 ), .A(
        \MCD/insdec_1/n4249 ), .B(\MCD/insdec_1/n4239 ) );
    snl_invx05 \MCD/insdec_1/U288  ( .ZN(\MCD/insdec_1/n4236 ), .A(
        \MCD/insdec_1/n4223 ) );
    snl_muxi21x1 \MCD/insdec_1/U318  ( .ZN(\MCD/insdec_1/n4210 ), .A(
        \MCD/insdec_1/n4203 ), .B(\MCD/insdec_1/n4233 ), .S(
        \MCD/insdec_1/n4244 ) );
    snl_invx05 \MCD/insdec_1/U242  ( .ZN(\MCD/insdec_1/n4185 ), .A(
        \stream4[46] ) );
    snl_muxi21x1 \MCD/insdec_1/U265  ( .ZN(\MCD/insdec_1/n4175 ), .A(
        \MCD/insdec_1/n4230 ), .B(\MCD/insdec_1/n4232 ), .S(\stream4[57] ) );
    snl_invx05 \MCD/insdec_1/U280  ( .ZN(\MCD/insdec_1/n4280 ), .A(
        \MCD/insdec_1/n4251 ) );
    snl_nand03x0 \MCD/insdec_1/U310  ( .ZN(\MCD/insdec_1/n4276 ), .A(
        \MCD/insdec_1/n4279 ), .B(\MCD/insdec_1/n4219 ), .C(
        \MCD/insdec_1/n4220 ) );
    snl_nor02x1 \MCD/insdec_1/U182  ( .ZN(baccsel), .A(\MCD/insdec_1/n4177 ), 
        .B(\MCD/insdec_1/n4178 ) );
    snl_nor03x0 \MCD/insdec_1/U185  ( .ZN(all0bsel), .A(\MCD/insdec_1/n4187 ), 
        .B(ph_saexe_sth), .C(\MCD/insdec_1/n4182 ) );
    snl_aoi033x0 \MCD/insdec_1/U202  ( .ZN(\MCD/insdec_1/n4176 ), .A(
        \MCD/insdec_1/n4224 ), .B(\MCD/insdec_1/n4225 ), .C(\stream4[51] ), 
        .D(\MCD/insdec_1/n4226 ), .E(\MCD/insdec_1/n4227 ), .F(\stream4[49] )
         );
    snl_muxi21x1 \MCD/insdec_1/U210  ( .ZN(\MCD/insdec_1/n4234 ), .A(
        \MCD/insdec_1/n4243 ), .B(\MCD/insdec_1/n4242 ), .S(
        \MCD/insdec_1/n4244 ) );
    snl_aoi022x1 \MCD/insdec_1/U259  ( .ZN(\MCD/insdec_1/n4260 ), .A(
        \MCD/insdec_1/n4228 ), .B(\stream4[33] ), .C(\MCD/insdec_1/n4271 ), 
        .D(\MCD/insdec_1/n4247 ) );
    snl_nand02x1 \MCD/insdec_1/U237  ( .ZN(\MCD/insdec_1/n4161 ), .A(
        \MCD/insdec_1/n4170 ), .B(\MCD/insdec_1/n4224 ) );
    snl_invx05 \MCD/insdec_1/U225  ( .ZN(\MCD/insdec_1/n4252 ), .A(stage_b) );
    snl_invx05 \MCD/insdec_1/U250  ( .ZN(\MCD/insdec_1/n4265 ), .A(
        \stream4[42] ) );
    snl_nand03x0 \MCD/insdec_1/U277  ( .ZN(\MCD/insdec_1/n4214 ), .A(
        \MCD/insdec_1/n4280 ), .B(\MCD/insdec_1/n4229 ), .C(stage_b) );
    snl_invx05 \MCD/insdec_1/U289  ( .ZN(\MCD/insdec_1/n4211 ), .A(
        \stream4[41] ) );
    snl_muxi21x1 \MCD/insdec_1/U319  ( .ZN(\MCD/insdec_1/n4275 ), .A(
        \MCD/insdec_1/n4273 ), .B(\MCD/insdec_1/n4213 ), .S(\stream4[47] ) );
    snl_invx05 \MCD/insdec_1/U219  ( .ZN(\MCD/insdec_1/n4239 ), .A(
        \stream4[32] ) );
    snl_invx05 \MCD/insdec_1/U292  ( .ZN(\MCD/insdec_1/n4237 ), .A(
        \MCD/insdec_1/n4263 ) );
    snl_oai012x1 \MCD/insdec_1/U302  ( .ZN(\MCD/insdec_1/n4164 ), .A(
        \stream4[39] ), .B(\stream4[37] ), .C(\MCD/insdec_1/n4170 ) );
    snl_invx05 \MCD/insdec_1/U295  ( .ZN(\MCD/insdec_1/n4259 ), .A(
        \MCD/insdec_1/n4254 ) );
    snl_invx05 \MCD/insdec_1/U305  ( .ZN(\poalufnc[1] ), .A(
        \MCD/insdec_1/n4169 ) );
    snl_invx05 \MCD/insdec_1/U239  ( .ZN(\MCD/insdec_1/n4166 ), .A(
        \stream4[37] ) );
    snl_invx05 \MCD/insdec_1/U322  ( .ZN(\MCD/insdec_1/n4282 ), .A(
        \stream4[36] ) );
    snl_nand14x0 \MCD/insdec_1/U175  ( .ZN(\poalufnc[3] ), .A(\stream4[38] ), 
        .B(\MCD/insdec_1/n4164 ), .C(\MCD/insdec_1/n4158 ), .D(
        \MCD/insdec_1/n4165 ) );
    snl_aoi012x1 \MCD/insdec_1/U199  ( .ZN(\MCD/insdec_1/n4221 ), .A(
        \MCD/insdec_1/n4222 ), .B(\MCD/insdec_1/n4223 ), .C(
        \MCD/insdec_1/n4202 ) );
    snl_nor02x1 \MCD/insdec_1/U205  ( .ZN(\MCD/insdec_1/n4232 ), .A(
        \MCD/insdec_1/n4233 ), .B(\MCD/insdec_1/n4234 ) );
    snl_invx05 \MCD/insdec_1/U222  ( .ZN(\MCD/insdec_1/n4250 ), .A(
        \MCD/insdec_1/ciff ) );
    snl_nor02x1 \MCD/insdec_1/U257  ( .ZN(\MCD/insdec_1/n4269 ), .A(
        \MCD/insdec_1/n4266 ), .B(\MCD/insdec_1/n4248 ) );
    snl_or04x1 \MCD/insdec_1/U270  ( .Z(\MCD/insdec_1/n4196 ), .A(
        \MCD/insdec_1/n4173 ), .B(\poalufnc[0] ), .C(\poalufnc[2] ), .D(
        \poalufnc[4] ) );
    snl_invx05 \MCD/insdec_1/U217  ( .ZN(\MCD/insdec_1/n4246 ), .A(
        \stream4[34] ) );
    snl_oa012x1 \MCD/insdec_1/U230  ( .Z(\MCD/insdec_1/n4216 ), .A(
        \MCD/insdec_1/n4200 ), .B(\MCD/insdec_1/n4255 ), .C(
        \MCD/insdec_1/n4257 ) );
    snl_invx05 \MCD/insdec_1/U279  ( .ZN(\MCD/insdec_1/n4172 ), .A(
        \MCD/insdec_1/n4207 ) );
    snl_nor02x1 \MCD/insdec_1/U190  ( .ZN(\MCD/insdec_1/n4198 ), .A(
        \stream4[55] ), .B(\MCD/insdec_1/n4199 ) );
    snl_invx05 \MCD/insdec_1/U245  ( .ZN(\MCD/insdec_1/n4227 ), .A(
        \stream4[48] ) );
    snl_oai013x0 \MCD/insdec_1/U262  ( .ZN(\MCD/insdec_1/n4195 ), .A(
        \MCD/insdec_1/n4182 ), .B(\stream4[44] ), .C(\MCD/insdec_1/n4274 ), 
        .D(\MCD/insdec_1/n4275 ) );
    snl_invx05 \MCD/insdec_1/U287  ( .ZN(eaccasel), .A(\MCD/insdec_1/n4186 )
         );
    snl_muxi21x1 \MCD/insdec_1/U317  ( .ZN(\MCD/insdec_1/n4271 ), .A(
        \stream4[32] ), .B(\MCD/insdec_1/n4270 ), .S(\MCD/insdec_1/bacc ) );
    snl_aoi022x1 \MCD/insdec_1/U207  ( .ZN(\MCD/insdec_1/n4238 ), .A(
        \MCD/insdec_1/ciff ), .B(\stream4[32] ), .C(pk_sign_h), .D(
        \MCD/insdec_1/n4239 ) );
    snl_nand12x1 \MCD/insdec_1/U220  ( .ZN(\MCD/insdec_1/n4248 ), .A(
        \stream4[59] ), .B(\stream4[58] ) );
    snl_or03x1 \MCD/insdec_1/U269  ( .Z(\MCD/insdec_1/n4277 ), .A(
        \poshtfnc[1] ), .B(\poshtfnc[2] ), .C(\poshtfnc[0] ) );
    snl_nand03x0 \MCD/insdec_1/U272  ( .ZN(\MCD/insdec_1/n4279 ), .A(
        \MCD/insdec_1/n4280 ), .B(\MCD/insdec_1/n4229 ), .C(
        \MCD/insdec_1/n4278 ) );
    snl_and02x2 \MCD/insdec_1/U170  ( .Z(eaccbsel), .A(\MCD/insdec_1/n4191 ), 
        .B(\MCD/insdec_1/n4165 ) );
    snl_nor03x0 \MCD/insdec_1/U177  ( .ZN(\MCD/insdec_1/n4169 ), .A(
        \MCD/insdec_1/n4170 ), .B(ph_saexe_sth), .C(\stream4[36] ) );
    snl_nor02x1 \MCD/insdec_1/U180  ( .ZN(ltffsel), .A(ph_saexe_sth), .B(
        \MCD/insdec_1/n4175 ) );
    snl_ao022x1 \MCD/insdec_1/U255  ( .Z(\MCD/insdec_1/n4266 ), .A(
        \MCD/insdec_1/n4238 ), .B(\MCD/insdec_1/n4246 ), .C(
        \MCD/insdec_1/n4267 ), .D(\stream4[34] ) );
    snl_aoi012x1 \MCD/insdec_1/U192  ( .ZN(\MCD/insdec_1/n4160 ), .A(
        \MCD/insdec_1/n4201 ), .B(\MCD/insdec_1/n4202 ), .C(
        \MCD/insdec_1/n4203 ) );
    snl_invx05 \MCD/insdec_1/U297  ( .ZN(\MCD/insdec_1/n4217 ), .A(
        \MCD/insdec_1/n4256 ) );
    snl_invx05 \MCD/insdec_1/U320  ( .ZN(\MCD/insdec_1/n4193 ), .A(
        \MCD/insdec_1/n4190 ) );
    snl_nor02x1 \MCD/insdec_1/U307  ( .ZN(\MCD/insdec_1/n4233 ), .A(
        \MCD/insdec_1/n4224 ), .B(\MCD/insdec_1/n4159 ) );
    snl_nor02x1 \MCD/insdec_1/U229  ( .ZN(\MCD/insdec_1/n4256 ), .A(
        \MCD/insdec_1/n4251 ), .B(\MCD/insdec_1/n4229 ) );
    snl_nor03x0 \MCD/insdec_1/U285  ( .ZN(wexacc), .A(\MCD/insdec_1/n4179 ), 
        .B(\MCD/insdec_1/n4190 ), .C(\MCD/insdec_1/n4180 ) );
    snl_aoi022x1 \MCD/insdec_1/U315  ( .ZN(\MCD/insdec_1/n4267 ), .A(
        \MCD/insdec_1/bacc ), .B(\MCD/insdec_1/n4239 ), .C(
        \MCD/insdec_1/n4250 ), .D(\stream4[32] ) );
    snl_mux21x1 \MCD/insdec_1/U260  ( .Z(\MCD/insdec_1/n4272 ), .A(
        \MCD/insdec_1/n4233 ), .B(\MCD/insdec_1/n4203 ), .S(
        \MCD/insdec_1/n4244 ) );
    snl_nor03x0 \MCD/insdec_1/U189  ( .ZN(srctype0), .A(\stream4[53] ), .B(
        \stream4[54] ), .C(\stream4[52] ) );
    snl_nor04x0 \MCD/insdec_1/U215  ( .ZN(\MCD/insdec_1/n4212 ), .A(
        \MCD/insdec_1/n4236 ), .B(\stream4[43] ), .C(\stream4[41] ), .D(
        \stream4[42] ) );
    snl_nand03x0 \MCD/insdec_1/U247  ( .ZN(\MCD/insdec_1/n4181 ), .A(
        \stream4[44] ), .B(\MCD/insdec_1/n4223 ), .C(\MCD/insdec_1/n4263 ) );
    snl_nor02x1 \MCD/insdec_1/U232  ( .ZN(\MCD/insdec_1/n4170 ), .A(
        \MCD/insdec_1/n4223 ), .B(ph_saexe_sth) );
    snl_invx05 \MCD/insdec_1/U212  ( .ZN(\MCD/insdec_1/n4199 ), .A(
        \stream4[56] ) );
    snl_invx05 \MCD/insdec_1/U235  ( .ZN(\MCD/insdec_1/n4171 ), .A(
        \stream4[35] ) );
    snl_nor02x1 \MCD/insdec_1/U240  ( .ZN(\MCD/insdec_1/n4207 ), .A(
        \MCD/insdec_1/n4236 ), .B(ph_saexe_sth) );
    snl_nand14x0 \MCD/insdec_1/U299  ( .ZN(\MCD/insdec_1/n4261 ), .A(
        \MCD/insdec_1/n4248 ), .B(\MCD/insdec_1/n4238 ), .C(
        \MCD/insdec_1/n4247 ), .D(\MCD/insdec_1/n4246 ) );
    snl_invx05 \MCD/insdec_1/U309  ( .ZN(\MCD/insdec_1/n4177 ), .A(
        \MCD/insdec_1/n4281 ) );
    snl_nand12x8 \MCD/insdec_1/U171  ( .ZN(po_arsel_h), .A(accasel), .B(
        \MCD/insdec_1/n4186 ) );
    snl_nor02x1 \MCD/insdec_1/U179  ( .ZN(ciffsel), .A(ph_saexe_sth), .B(
        \MCD/insdec_1/n4174 ) );
    snl_oa012x1 \MCD/insdec_1/U187  ( .Z(po_reacl_h), .A(\MCD/insdec_1/n4191 ), 
        .B(\MCD/insdec_1/n4192 ), .C(\MCD/insdec_1/n4193 ) );
    snl_nor02x1 \MCD/insdec_1/U195  ( .ZN(\MCD/insdec_1/n4208 ), .A(
        \poalufnc[4] ), .B(\MCD/insdec_1/n4194 ) );
    snl_aoi022x1 \MCD/insdec_1/U267  ( .ZN(\MCD/insdec_1/n4187 ), .A(
        \MCD/insdec_1/n4276 ), .B(\stream4[44] ), .C(\MCD/insdec_1/n4235 ), 
        .D(\MCD/insdec_1/n4241 ) );
    snl_and23x0 \MCD/insdec_1/U282  ( .Z(srctype2), .A(\stream4[52] ), .B(
        \stream4[54] ), .C(\stream4[53] ) );
    snl_nand12x1 \MCD/insdec_1/U312  ( .ZN(\MCD/insdec_1/n4189 ), .A(
        \MCD/insdec_1/n4184 ), .B(\MCD/insdec_1/n4263 ) );
    snl_muxi21x1 \MCD/insdec_1/U209  ( .ZN(\MCD/insdec_1/n4231 ), .A(
        \MCD/insdec_1/n4242 ), .B(\MCD/insdec_1/n4243 ), .S(
        \MCD/insdec_1/n4244 ) );
    snl_ao1b1b2x0 \MCD/insdec_1/U290  ( .Z(\MCD/insdec_1/n4168 ), .A(
        \MCD/insdec_1/n4204 ), .B(\MCD/insdec_1/n4203 ), .C(
        \MCD/insdec_1/n4214 ), .D(\MCD/insdec_1/n4158 ) );
    snl_invx05 \MCD/insdec_1/U300  ( .ZN(\MCD/insdec_1/n4205 ), .A(
        \MCD/insdec_1/n4202 ) );
    snl_nor02x1 \MCD/insdec_1/U252  ( .ZN(\MCD/insdec_1/n4191 ), .A(
        \MCD/insdec_1/n4181 ), .B(\stream4[45] ) );
    snl_nor02x1 \MCD/insdec_1/U275  ( .ZN(\poshtfnc[0] ), .A(
        \MCD/insdec_1/n4239 ), .B(\MCD/insdec_1/n4236 ) );
    snl_nor02x1 \MCD/insdec_1/U194  ( .ZN(\MCD/insdec_1/n4162 ), .A(
        \MCD/insdec_1/n4206 ), .B(\MCD/insdec_1/n4207 ) );
    snl_nor02x1 \MCD/insdec_1/U200  ( .ZN(\MCD/insdec_1/n4197 ), .A(wexacc), 
        .B(wacc) );
    snl_nor02x1 \MCD/insdec_1/U227  ( .ZN(\MCD/insdec_1/n4254 ), .A(
        \MCD/insdec_1/n4248 ), .B(\MCD/insdec_1/n4246 ) );
    snl_nor03x0 \MCD/insdec_1/U249  ( .ZN(\MCD/insdec_1/n4194 ), .A(
        \poalufnc[1] ), .B(\poalufnc[2] ), .C(\poalufnc[0] ) );
    snl_nor02x1 \MCD/insdec_1/U283  ( .ZN(accasel), .A(\MCD/insdec_1/n4188 ), 
        .B(ph_saexe_sth) );
    snl_oai012x1 \MCD/insdec_1/U313  ( .ZN(\MCD/insdec_1/n4226 ), .A(
        \MCD/insdec_1/n4236 ), .B(\MCD/insdec_1/n4264 ), .C(
        \MCD/insdec_1/n4205 ) );
    snl_aoi022x1 \MCD/insdec_1/U208  ( .ZN(\MCD/insdec_1/n4240 ), .A(
        \stream4[44] ), .B(\MCD/insdec_1/n4182 ), .C(\MCD/insdec_1/n4241 ), 
        .D(\stream4[45] ) );
    snl_invx05 \MCD/insdec_1/U241  ( .ZN(\MCD/insdec_1/n4182 ), .A(
        \stream4[45] ) );
    snl_aoi1b12x0 \MCD/insdec_1/U178  ( .ZN(po_cmfsel_h), .A(\poalufnc[2] ), 
        .B(\poalufnc[1] ), .C(\poalufnc[4] ), .D(\MCD/insdec_1/n4173 ) );
    snl_aoi033x0 \MCD/insdec_1/U201  ( .ZN(\MCD/insdec_1/n4183 ), .A(
        \stream4[48] ), .B(\MCD/insdec_1/n4202 ), .C(\stream4[49] ), .D(
        \stream4[50] ), .E(\MCD/insdec_1/n4224 ), .F(\stream4[51] ) );
    snl_invx05 \MCD/insdec_1/U213  ( .ZN(\MCD/insdec_1/n4245 ), .A(
        \stream4[55] ) );
    snl_oa122x1 \MCD/insdec_1/U234  ( .Z(\MCD/insdec_1/n4220 ), .A(
        \MCD/insdec_1/n4255 ), .B(\MCD/insdec_1/n4258 ), .C(
        \MCD/insdec_1/n4259 ), .D(\MCD/insdec_1/n4260 ), .E(
        \MCD/insdec_1/n4261 ) );
    snl_muxi21x1 \MCD/insdec_1/U266  ( .ZN(\MCD/insdec_1/n4174 ), .A(
        \MCD/insdec_1/n4232 ), .B(\MCD/insdec_1/n4230 ), .S(\stream4[57] ) );
    snl_and02x1 \MCD/insdec_1/U226  ( .Z(\MCD/insdec_1/n4253 ), .A(
        \MCD/insdec_1/n4249 ), .B(\MCD/insdec_1/n4251 ) );
    snl_invx05 \MCD/insdec_1/U298  ( .ZN(\MCD/insdec_1/n4262 ), .A(
        \MCD/insdec_1/n4224 ) );
    snl_oai023x0 \MCD/insdec_1/U308  ( .ZN(\MCD/insdec_1/n4281 ), .A(
        \MCD/insdec_1/n4272 ), .B(\stream4[42] ), .C(\stream4[43] ), .D(
        \stream4[40] ), .E(\MCD/insdec_1/n4209 ) );
    snl_ffqrnx1 \MCD/insdec_1/bacc_reg  ( .Q(\MCD/insdec_1/bacc ), .D(pk_bacch
        ), .RN(n10733), .CP(SCLK) );
    snl_oa023x1 \MCD/insdec_1/U248  ( .Z(\MCD/insdec_1/n4188 ), .A(
        \MCD/insdec_1/n4221 ), .B(\stream4[49] ), .C(\stream4[48] ), .D(
        \MCD/insdec_1/n4262 ), .E(\MCD/insdec_1/n4264 ) );
    snl_nor04x0 \MCD/insdec_1/U253  ( .ZN(\MCD/insdec_1/n4192 ), .A(
        \MCD/insdec_1/n4227 ), .B(\MCD/insdec_1/n4264 ), .C(
        \MCD/insdec_1/n4236 ), .D(\stream4[49] ) );
    snl_oai122x2 \MCD/insdec_1/U164  ( .ZN(\poalufnc[0] ), .A(
        \MCD/insdec_1/n4167 ), .B(\MCD/insdec_1/n4161 ), .C(
        \MCD/insdec_1/n4171 ), .D(\MCD/insdec_1/n4172 ), .E(
        \MCD/insdec_1/n4168 ) );
    snl_nor02x1 \MCD/insdec_1/U181  ( .ZN(all0asel), .A(ph_saexe_sth), .B(
        \MCD/insdec_1/n4176 ) );
    snl_aoi012x1 \MCD/insdec_1/U186  ( .ZN(po_raccl_h), .A(
        \MCD/insdec_1/n4188 ), .B(\MCD/insdec_1/n4189 ), .C(
        \MCD/insdec_1/n4190 ) );
    snl_nor02x1 \MCD/insdec_1/U274  ( .ZN(\poshtfnc[1] ), .A(
        \MCD/insdec_1/n4247 ), .B(\MCD/insdec_1/n4236 ) );
    snl_invx05 \MCD/insdec_1/U291  ( .ZN(\MCD/insdec_1/n4179 ), .A(
        \MCD/insdec_1/n4212 ) );
    snl_and02x1 \MCD/insdec_1/U301  ( .Z(\MCD/insdec_1/n4203 ), .A(
        \MCD/insdec_1/n4205 ), .B(\MCD/insdec_1/n4279 ) );
    snl_nor02x1 \MCD/insdec_1/U273  ( .ZN(\poshtfnc[2] ), .A(
        \MCD/insdec_1/n4246 ), .B(\MCD/insdec_1/n4236 ) );
    snl_invx05 \MCD/insdec_1/U296  ( .ZN(\MCD/insdec_1/n4278 ), .A(
        \MCD/insdec_1/n4218 ) );
    snl_oa012x1 \MCD/insdec_1/U306  ( .Z(\MCD/insdec_1/n4244 ), .A(srctype1), 
        .B(srctype2), .C(\MCD/insdec_1/n4256 ) );
    snl_invx05 \MCD/insdec_1/U321  ( .ZN(\MCD/insdec_1/n4241 ), .A(
        \stream4[44] ) );
    snl_oai122x0 \MCD/insdec_1/U176  ( .ZN(\poalufnc[2] ), .A(
        \MCD/insdec_1/n4162 ), .B(\MCD/insdec_1/n4166 ), .C(
        \MCD/insdec_1/n4167 ), .D(\MCD/insdec_1/n4161 ), .E(
        \MCD/insdec_1/n4168 ) );
    snl_and23x0 \MCD/insdec_1/U188  ( .Z(po_opcsel_h), .A(\poalufnc[4] ), .B(
        \MCD/insdec_1/n4173 ), .C(\MCD/insdec_1/n4194 ) );
    snl_nor02x1 \MCD/insdec_1/U206  ( .ZN(\MCD/insdec_1/n4235 ), .A(
        \MCD/insdec_1/n4236 ), .B(\MCD/insdec_1/n4237 ) );
    snl_invx05 \MCD/insdec_1/U254  ( .ZN(\MCD/insdec_1/n4225 ), .A(
        \stream4[50] ) );
    snl_ao022x1 \MCD/insdec_1/U268  ( .Z(\MCD/insdec_1/n4258 ), .A(
        \MCD/insdec_1/ciff ), .B(\MCD/insdec_1/bacc ), .C(\pk_stat_h[18] ), 
        .D(ph_piosl_h) );
    snl_oai012x1 \MCD/insdec_1/U214  ( .ZN(\MCD/insdec_1/n4190 ), .A(
        \MCD/insdec_1/n4198 ), .B(exetype1), .C(\MCD/insdec_1/n4165 ) );
    snl_nor03x0 \MCD/insdec_1/U221  ( .ZN(\MCD/insdec_1/n4249 ), .A(
        \MCD/insdec_1/n4247 ), .B(\stream4[34] ), .C(\MCD/insdec_1/n4248 ) );
    snl_nand02x1 \MCD/insdec_1/U233  ( .ZN(\MCD/insdec_1/n4218 ), .A(stage_2), 
        .B(\MCD/insdec_1/n4252 ) );
    snl_nor03x0 \MCD/insdec_1/U261  ( .ZN(\MCD/insdec_1/n4273 ), .A(
        \MCD/insdec_1/n4185 ), .B(\MCD/insdec_1/n4240 ), .C(
        \MCD/insdec_1/n4236 ) );
    snl_aoi012x1 \MCD/insdec_1/U193  ( .ZN(\MCD/insdec_1/n4204 ), .A(
        \stream4[36] ), .B(\MCD/insdec_1/n4171 ), .C(\MCD/insdec_1/n4205 ) );
    snl_nor02x1 \MCD/insdec_1/U246  ( .ZN(\MCD/insdec_1/n4263 ), .A(
        \stream4[46] ), .B(\stream4[47] ) );
    snl_nand03x0 \MCD/insdec_1/U228  ( .ZN(\MCD/insdec_1/n4255 ), .A(
        \stream4[32] ), .B(\stream4[33] ), .C(\MCD/insdec_1/n4254 ) );
    snl_oa113x1 \MCD/insdec_1/U284  ( .Z(wacc), .A(\MCD/insdec_1/n4277 ), .B(
        \MCD/insdec_1/n4173 ), .C(\MCD/insdec_1/n4208 ), .D(
        \MCD/insdec_1/n4193 ), .E(\MCD/insdec_1/n4281 ) );
    snl_aoi022x1 \MCD/insdec_1/U314  ( .ZN(\MCD/insdec_1/n4201 ), .A(
        \stream4[35] ), .B(\MCD/insdec_1/n4282 ), .C(\MCD/insdec_1/n4171 ), 
        .D(\stream4[36] ) );
    snl_oai112x0 \MAIN/MCD/U55  ( .ZN(\MAIN/MCD/nst[0] ), .A(\MAIN/MCD/dst[1] 
        ), .B(\MAIN/MCD/n3367 ), .C(\MAIN/MCD/n3368 ), .D(\MAIN/MCD/n3369 ) );
    snl_nor02x1 \MAIN/MCD/U61  ( .ZN(\MAIN/MCD/n3367 ), .A(\MAIN/st_decctl ), 
        .B(\MAIN/MCD/n3381 ) );
    snl_invx05 \MAIN/MCD/U68  ( .ZN(\MAIN/MCD/n3378 ), .A(\MAIN/MCD/dst[0] )
         );
    snl_muxi21x1 \MAIN/MCD/U73  ( .ZN(\MAIN/MCD/n3387 ), .A(\MAIN/MCD/n3388 ), 
        .B(\MAIN/MCD/n3389 ), .S(po_sprtrs_h) );
    snl_nand12x1 \MAIN/MCD/U84  ( .ZN(\MAIN/MCD/n3388 ), .A(po_oprtrs_h), .B(
        \MAIN/cstregw_inhibith ) );
    snl_nor02x1 \MAIN/MCD/U66  ( .ZN(\MAIN/MCD/n3383 ), .A(\MAIN/MCD/n3373 ), 
        .B(\MAIN/EXCEP_EXT ) );
    snl_nand02x1 \MAIN/MCD/U67  ( .ZN(\MAIN/MCD/n3371 ), .A(\MAIN/MCD/dst[1] ), 
        .B(\MAIN/MCD/n3378 ) );
    snl_muxi21x1 \MAIN/MCD/U74  ( .ZN(\MAIN/MCD/n3390 ), .A(\MAIN/MCD/n3380 ), 
        .B(\MAIN/MCD/n3391 ), .S(po_sprtrs_h) );
    snl_invx05 \MAIN/MCD/U83  ( .ZN(\MAIN/MCD/n3397 ), .A(\MAIN/MCD/n3371 ) );
    snl_aoi022x1 \MAIN/MCD/U91  ( .ZN(\MAIN/MCD/n3379 ), .A(\MAIN/MCD/n3393 ), 
        .B(\MAIN/MCD/dst[2] ), .C(\MAIN/MCD/n3395 ), .D(\MAIN/MCD/n3374 ) );
    snl_ffqrnx1 \MAIN/MCD/dst_reg[1]  ( .Q(\MAIN/MCD/dst[1] ), .D(
        \MAIN/MCD/nst[1] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \MAIN/MCD/U82  ( .ZN(\MAIN/MCD/n3384 ), .A(\MAIN/MCD/n3377 ) );
    snl_aoi022x1 \MAIN/MCD/U69  ( .ZN(\MAIN/MCD/n3368 ), .A(\MAIN/MCD/n3378 ), 
        .B(\MAIN/MCD/dst[2] ), .C(\MAIN/MCD/n3376 ), .D(\MAIN/MCD/n3384 ) );
    snl_nor02x1 \MAIN/MCD/U75  ( .ZN(\MAIN/MCD/n3392 ), .A(
        \MAIN/dprw_inhibith ), .B(\MAIN/MCD/n3387 ) );
    snl_muxi21x1 \MAIN/MCD/U90  ( .ZN(\MAIN/MCD/n3398 ), .A(\MAIN/MCD/n3390 ), 
        .B(\MAIN/MCD/n3392 ), .S(po_dprtrs_h) );
    snl_nand12x1 \MAIN/MCD/U72  ( .ZN(\MAIN/MCD/n3385 ), .A(\MAIN/EXCEP_EXT ), 
        .B(\MAIN/MCD/n3386 ) );
    snl_oai012x1 \MAIN/MCD/U56  ( .ZN(\MAIN/MCD/nst[1] ), .A(\MAIN/MCD/dst[2] 
        ), .B(\MAIN/MCD/n3370 ), .C(\MAIN/MCD/n3368 ) );
    snl_oai133x0 \MAIN/MCD/U57  ( .ZN(\MAIN/MCD/nst[2] ), .A(\MAIN/MCD/n3371 ), 
        .B(\MAIN/MCD/n3372 ), .C(\MAIN/MCD/n3373 ), .D(\MAIN/MCD/n3374 ), .E(
        \MAIN/MCD/dst[1] ), .F(\MAIN/MCD/n3375 ), .G(\MAIN/MCD/n3368 ) );
    snl_oa012x1 \MAIN/MCD/U60  ( .Z(\MAIN/MCD/n3380 ), .A(
        \MAIN/cstregw_inhibith ), .B(\MAIN/astregw_inhibith ), .C(po_oprtrs_h)
         );
    snl_nand12x1 \MAIN/MCD/U85  ( .ZN(\MAIN/MCD/n3396 ), .A(\MAIN/st_decctl ), 
        .B(\MAIN/MCD/n3386 ) );
    snl_oai013x0 \MAIN/MCD/U58  ( .ZN(\MAIN/dec_end ), .A(\MAIN/MCD/n3376 ), 
        .B(\MAIN/MCD/n3377 ), .C(\MAIN/MCD/n3378 ), .D(\MAIN/MCD/n3379 ) );
    snl_or02x1 \MAIN/MCD/U59  ( .Z(\MAIN/MCD/stage_a154 ), .A(
        \MAIN/MCD/nst[1] ), .B(\MAIN/MCD/nst[0] ) );
    snl_aoi012x1 \MAIN/MCD/U62  ( .ZN(\MAIN/MCD/n3370 ), .A(\MAIN/MCD/dst[1] ), 
        .B(\MAIN/MCD/n3382 ), .C(\MAIN/MCD/dst[0] ) );
    snl_invx05 \MAIN/MCD/U70  ( .ZN(\MAIN/MCD/n3376 ), .A(\MAIN/POL_STH ) );
    snl_aoi023x0 \MAIN/MCD/U79  ( .ZN(\MAIN/MCD/n3369 ), .A(\MAIN/MCD/n3383 ), 
        .B(\MAIN/MCD/n3396 ), .C(\MAIN/MCD/n3397 ), .D(\MAIN/st_decctl ), .E(
        \MAIN/MCD/n3384 ) );
    snl_invx05 \MAIN/MCD/U87  ( .ZN(\MAIN/MCD/n3382 ), .A(\MAIN/MCD/n3383 ) );
    snl_invx05 \MAIN/MCD/U65  ( .ZN(\MAIN/MCD/n3373 ), .A(\MAIN/decend_en ) );
    snl_invx05 \MAIN/MCD/U80  ( .ZN(\MAIN/MCD/n3389 ), .A(\MAIN/sprw_inhibith 
        ) );
    snl_nor02x1 \MAIN/MCD/U77  ( .ZN(\MAIN/MCD/n3393 ), .A(\MAIN/MCD/dst[1] ), 
        .B(\MAIN/MCD/n3394 ) );
    snl_nand02x1 \MAIN/MCD/U89  ( .ZN(\MAIN/MCD/n3391 ), .A(\MAIN/MCD/n3388 ), 
        .B(\MAIN/MCD/n3389 ) );
    snl_nand14x0 \MAIN/MCD/U64  ( .ZN(\MAIN/MCD/n3377 ), .A(\MAIN/WP_PC ), .B(
        pk_pexe01_h), .C(\MAIN/MCD/dst[1] ), .D(\MAIN/MCD/dst[2] ) );
    snl_nand12x1 \MAIN/MCD/U81  ( .ZN(\MAIN/MCD/n3386 ), .A(po_mode01_h), .B(
        \MAIN/MCD/n3398 ) );
    snl_ffqrnx1 \MAIN/MCD/dst_reg[0]  ( .Q(\MAIN/MCD/dst[0] ), .D(
        \MAIN/MCD/nst[0] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_ffqrnx1 \MAIN/MCD/stage_a_reg  ( .Q(stage_a), .D(\MAIN/MCD/stage_a154 
        ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_aoi022x1 \MAIN/MCD/U76  ( .ZN(\MAIN/MCD/n3381 ), .A(\MAIN/MCD/n3375 ), 
        .B(\MAIN/MCD/dst[2] ), .C(\MAIN/MCD/n3378 ), .D(\MAIN/MCD/n3374 ) );
    snl_invx05 \MAIN/MCD/U88  ( .ZN(\MAIN/MCD/n3372 ), .A(\MAIN/MCD/n3385 ) );
    snl_invx05 \MAIN/MCD/U63  ( .ZN(\MAIN/MCD/n3374 ), .A(\MAIN/MCD/dst[2] )
         );
    snl_nor04x0 \MAIN/MCD/U71  ( .ZN(\MAIN/MCD/n3375 ), .A(
        \MAIN/cstregw_inhibith ), .B(\MAIN/astregw_inhibith ), .C(
        \MAIN/sprw_inhibith ), .D(\MAIN/dprw_inhibith ) );
    snl_nor03x0 \MAIN/MCD/U78  ( .ZN(\MAIN/MCD/n3395 ), .A(\MAIN/MCD/n3385 ), 
        .B(\MAIN/MCD/n3373 ), .C(\MAIN/MCD/n3371 ) );
    snl_invx05 \MAIN/MCD/U86  ( .ZN(\MAIN/MCD/n3394 ), .A(\MAIN/MCD/n3375 ) );
    snl_ffqrnx1 \MAIN/MCD/dst_reg[2]  ( .Q(\MAIN/MCD/dst[2] ), .D(
        \MAIN/MCD/nst[2] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_bufx1 \REGF/pbmemcnt1/U206  ( .Z(\REGF/pbmemcnt1/n6441 ), .A(
        \REGF/n8052 ) );
    snl_and23x1 \REGF/pbmemcnt1/U207  ( .Z(\REGF/pbmemcnt1/n6443 ), .A(
        ph_schvx_h), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/n6447 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U210  ( .Z(\REGF/pbmemcnt1/upcnt_data392[9] ), 
        .A(\pk_stdat[9] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[9] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U211  ( .Z(\REGF/pbmemcnt1/upcnt_data392[8] ), 
        .A(\pk_stdat[8] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[8] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U216  ( .Z(\REGF/pbmemcnt1/upcnt_data392[3] ), 
        .A(\pk_stdat[3] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[3] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_oai012x1 \REGF/pbmemcnt1/U223  ( .ZN(\REGF/pbmemcnt1/n401 ), .A(
        \REGF/pbmemcnt1/end_flag ), .B(\REGF/pbmemcnt1/n6495 ), .C(
        \REGF/pbmemcnt1/n6446 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U231  ( .Z(\REGF/pbmemcnt1/down_data404[5] ), 
        .A(PDLIN[5]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[5] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_nand02x1 \REGF/pbmemcnt1/U238  ( .ZN(\REGF/pbmemcnt1/n6449 ), .A(
        \REGF/pbmemcnt1/n6453 ), .B(\REGF/pbmemcnt1/upcnt_data[2] ) );
    snl_sffqensnx2 \REGF/pbmemcnt1/end_flag_reg  ( .Q(
        \REGF/pbmemcnt1/end_flag ), .D(1'b1), .EN(\REGF/pbmemcnt1/n6495 ), 
        .SN(\REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/n6494 ), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_invx05 \REGF/pbmemcnt1/U244  ( .ZN(\REGF/pbmemcnt1/n6494 ), .A(
        \REGF/pbmemcnt1/n6444 ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[5]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[5] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[5] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[8]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[8] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[8] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[1]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[1] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[1] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemcnt1/U218  ( .Z(\REGF/pbmemcnt1/upcnt_data392[1] ), 
        .A(\pk_stdat[1] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[1] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U236  ( .Z(\REGF/pbmemcnt1/down_data404[0] ), 
        .A(PDLIN[0]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[0] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_or08x1 \REGF/pbmemcnt1/U243  ( .Z(\REGF/pbmemcnt1/n6444 ), .A(PDLIN[1]
        ), .B(PDLIN[0]), .C(PDLIN[3]), .D(PDLIN[2]), .E(PDLIN[5]), .F(PDLIN[4]
        ), .G(PDLIN[7]), .H(PDLIN[6]) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[3]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[3] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[3] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[11]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[11] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[11] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[7]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[7] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[7] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_oai013x0 \REGF/pbmemcnt1/U224  ( .ZN(\REGF/pbmemcnt1/n405[0] ), .A(
        \REGF/pbmemcnt1/n6447 ), .B(\REGF/pbmemcnt1/end_flag ), .C(
        \REGF/pbmemcnt1/n6448 ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_invx05 \REGF/pbmemcnt1/U242  ( .ZN(\REGF/pbmemcnt1/n6445 ), .A(
        \REGF/pbmemcnt1/n6495 ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[3]  ( .Q(
        \REGF/pbmemcnt1/down_data[3] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[3] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemcnt1/U217  ( .Z(\REGF/pbmemcnt1/upcnt_data392[2] ), 
        .A(\pk_stdat[2] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[2] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U219  ( .Z(\REGF/pbmemcnt1/upcnt_data392[0] ), 
        .A(\pk_stdat[0] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[0] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_or08x1 \REGF/pbmemcnt1/U225  ( .Z(\REGF/pbmemcnt1/n6447 ), .A(
        \REGF/pbmemcnt1/upcnt_data[5] ), .B(\REGF/pbmemcnt1/upcnt_data[4] ), 
        .C(\REGF/pbmemcnt1/upcnt_data[3] ), .D(\REGF/pbmemcnt1/upcnt_data[9] ), 
        .E(\REGF/pbmemcnt1/upcnt_data[7] ), .F(\REGF/pbmemcnt1/upcnt_data[6] ), 
        .G(\REGF/pbmemcnt1/n6449 ), .H(\REGF/pbmemcnt1/n6450 ) );
    snl_nor02x1 \REGF/pbmemcnt1/U237  ( .ZN(\REGF/pbmemcnt1/n6453 ), .A(
        \REGF/pbmemcnt1/upcnt_data[1] ), .B(\REGF/pbmemcnt1/upcnt_data[0] ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[7]  ( .Q(
        \REGF/pbmemcnt1/down_data[7] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[7] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_nand12x1 \REGF/pbmemcnt1/U222  ( .ZN(\REGF/pbmemcnt1/n6495 ), .A(
        \REGF/pbmemcnt1/n6447 ), .B(\REGF/pbmemcnt1/n6448 ) );
    snl_nand03x0 \REGF/pbmemcnt1/U239  ( .ZN(\REGF/pbmemcnt1/n6450 ), .A(
        \REGF/pbmemcnt1/upcnt_data[10] ), .B(\REGF/pbmemcnt1/upcnt_data[8] ), 
        .C(\REGF/pbmemcnt1/upcnt_data[11] ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[5]  ( .Q(
        \REGF/pbmemcnt1/down_data[5] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[5] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/time_delay_reg  ( .Q(\REGF/pk_sctio_h ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemcnt1/n6441 ), .SD(
        \REGF/pbmemcnt1/time_delay400 ), .SE(\REGF/pbmemcnt1/n401 ), .CP(SCLK)
         );
    snl_ao022x1 \REGF/pbmemcnt1/U230  ( .Z(\REGF/pbmemcnt1/down_data404[6] ), 
        .A(PDLIN[6]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[6] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[1]  ( .Q(
        \REGF/pbmemcnt1/down_data[1] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[1] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[0]  ( .Q(
        \REGF/pbmemcnt1/down_data[0] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[0] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemcnt1/U208  ( .Z(\REGF/pbmemcnt1/upcnt_data392[11] ), 
        .A(\pk_stdat[11] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[11] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U209  ( .Z(\REGF/pbmemcnt1/upcnt_data392[10] ), 
        .A(\pk_stdat[10] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[10] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U212  ( .Z(\REGF/pbmemcnt1/upcnt_data392[7] ), 
        .A(\pk_stdat[7] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[7] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U215  ( .Z(\REGF/pbmemcnt1/upcnt_data392[4] ), 
        .A(\pk_stdat[4] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[4] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_nand02x1 \REGF/pbmemcnt1/U220  ( .ZN(\REGF/pbmemcnt1/time_delay400 ), 
        .A(\pk_rwrit_h[2] ), .B(\REGF/pbmemcnt1/n6444 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U229  ( .Z(\REGF/pbmemcnt1/down_data404[7] ), 
        .A(PDLIN[7]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[7] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[4]  ( .Q(
        \REGF/pbmemcnt1/down_data[4] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[4] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemcnt1/U232  ( .Z(\REGF/pbmemcnt1/down_data404[4] ), 
        .A(PDLIN[4]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[4] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U235  ( .Z(\REGF/pbmemcnt1/down_data404[1] ), 
        .A(PDLIN[1]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[1] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_nor04x0 \REGF/pbmemcnt1/U240  ( .ZN(\REGF/pbmemcnt1/n6452 ), .A(
        \REGF/pbmemcnt1/down_data[7] ), .B(\REGF/pbmemcnt1/down_data[6] ), .C(
        \REGF/pbmemcnt1/down_data[5] ), .D(\REGF/pbmemcnt1/down_data[4] ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[6]  ( .Q(
        \REGF/pbmemcnt1/down_data[6] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[6] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_and03x1 \REGF/pbmemcnt1/U227  ( .Z(\REGF/pbmemcnt1/n6442 ), .A(
        \REGF/pbmemcnt1/n6447 ), .B(\REGF/pbmemcnt1/n6446 ), .C(ph_schvx_h) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/down_data_reg[2]  ( .Q(
        \REGF/pbmemcnt1/down_data[2] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/down_data404[2] ), .SE(
        \REGF/pbmemcnt1/n405[0] ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemcnt1/U213  ( .Z(\REGF/pbmemcnt1/upcnt_data392[6] ), 
        .A(\pk_stdat[6] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[6] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_ao022x1 \REGF/pbmemcnt1/U234  ( .Z(\REGF/pbmemcnt1/down_data404[2] ), 
        .A(PDLIN[2]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[2] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_and34x0 \REGF/pbmemcnt1/U241  ( .Z(\REGF/pbmemcnt1/n6451 ), .A(
        \REGF/pbmemcnt1/down_data[3] ), .B(\REGF/pbmemcnt1/down_data[2] ), .C(
        \REGF/pbmemcnt1/down_data[1] ), .D(\REGF/pbmemcnt1/down_data[0] ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[6]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[6] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[6] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_and02x1 \REGF/pbmemcnt1/U226  ( .Z(\REGF/pbmemcnt1/n6448 ), .A(
        \REGF/pbmemcnt1/n6451 ), .B(\REGF/pbmemcnt1/n6452 ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[10]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[10] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[10] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[2]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[2] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[2] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[9]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[9] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[9] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[0]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[0] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[0] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemcnt1/U214  ( .Z(\REGF/pbmemcnt1/upcnt_data392[5] ), 
        .A(\pk_stdat[5] ), .B(\REGF/pbmemcnt1/n6442 ), .C(
        \REGF/pbmemcnt1/upcnt_data283[5] ), .D(\REGF/pbmemcnt1/n6443 ) );
    snl_oai012x1 \REGF/pbmemcnt1/U221  ( .ZN(\REGF/pbmemcnt1/n393[0] ), .A(
        \REGF/pbmemcnt1/end_flag ), .B(\REGF/pbmemcnt1/n6445 ), .C(
        \REGF/pbmemcnt1/n6446 ) );
    snl_invx05 \REGF/pbmemcnt1/U228  ( .ZN(\REGF/pbmemcnt1/n6446 ), .A(
        \pk_rwrit_h[2] ) );
    snl_ao022x1 \REGF/pbmemcnt1/U233  ( .Z(\REGF/pbmemcnt1/down_data404[3] ), 
        .A(PDLIN[3]), .B(\pk_rwrit_h[2] ), .C(\REGF/pbmemcnt1/down_data274[3] 
        ), .D(\REGF/pbmemcnt1/n6446 ) );
    snl_sffqenrnx1 \REGF/pbmemcnt1/upcnt_data_reg[4]  ( .Q(
        \REGF/pbmemcnt1/upcnt_data[4] ), .D(1'b0), .EN(1'b1), .RN(
        \REGF/pbmemcnt1/n6441 ), .SD(\REGF/pbmemcnt1/upcnt_data392[4] ), .SE(
        \REGF/pbmemcnt1/n393[0] ), .CP(SCLK) );
    snl_and02x1 \SAEXE/SRCWT/U26  ( .Z(\SAEXE/SRCWT/nwst[1] ), .A(ph_lbend), 
        .B(\SAEXE/SRCWT/ewst[0] ) );
    snl_and23x0 \SAEXE/SRCWT/U28  ( .Z(\SAEXE/sa_start2 ), .A(
        \SAEXE/SRCWT/ewst[0] ), .B(\SAEXE/exec_end2 ), .C(\SAEXE/srcwt_st ) );
    snl_ffqrnx1 \SAEXE/SRCWT/ewst_reg[1]  ( .Q(\SAEXE/exec_end2 ), .D(
        \SAEXE/SRCWT/nwst[1] ), .RN(n10735), .CP(SCLK) );
    snl_ao012x1 \SAEXE/SRCWT/U27  ( .Z(\SAEXE/SRCWT/nwst[0] ), .A(
        \SAEXE/SRCWT/n85 ), .B(\SAEXE/SRCWT/ewst[0] ), .C(\SAEXE/sa_start2 )
         );
    snl_invx05 \SAEXE/SRCWT/U29  ( .ZN(\SAEXE/SRCWT/n85 ), .A(ph_lbend) );
    snl_ffqrnx1 \SAEXE/SRCWT/ewst_reg[0]  ( .Q(\SAEXE/SRCWT/ewst[0] ), .D(
        \SAEXE/SRCWT/nwst[0] ), .RN(n10735), .CP(SCLK) );
    snl_nor04x0 \MCD/adsel_1/U70  ( .ZN(po_raccen_h), .A(\MCD/adsel_1/n4283 ), 
        .B(\MCD/adsel_1/n4284 ), .C(\stream3[56] ), .D(\MCD/adsel_1/n4285 ) );
    snl_nor02x1 \MCD/adsel_1/U72  ( .ZN(wdpr), .A(\stream3[40] ), .B(
        \MCD/adsel_1/n4287 ) );
    snl_nor02x1 \MCD/adsel_1/U73  ( .ZN(wspr), .A(\MCD/adsel_1/n4287 ), .B(
        \MCD/adsel_1/n4288 ) );
    snl_nand02x1 \MCD/adsel_1/U74  ( .ZN(po_atchk_h), .A(\MCD/adsel_1/n4289 ), 
        .B(\MCD/adsel_1/n4290 ) );
    snl_aoi022x1 \MCD/adsel_1/U83  ( .ZN(\MCD/adsel_1/n4293 ), .A(
        \MCD/adsel_1/n4305 ), .B(\stream3[40] ), .C(\MCD/adsel_1/n4306 ), .D(
        \stream3[42] ) );
    snl_nor02x1 \MCD/adsel_1/U84  ( .ZN(\MCD/adsel_1/n4307 ), .A(
        \MCD/adsel_1/n4308 ), .B(\MCD/adsel_1/n4309 ) );
    snl_and34x0 \MCD/adsel_1/U96  ( .Z(po_ptrsel_h), .A(\MCD/adsel_1/n4332 ), 
        .B(\stream3[43] ), .C(\stream3[41] ), .D(po_mode01_h) );
    snl_nand02x1 \MCD/adsel_1/U113  ( .ZN(\MCD/adsel_1/n4343 ), .A(
        \MCD/adsel_1/n4337 ), .B(\MCD/adsel_1/n4344 ) );
    snl_nor02x1 \MCD/adsel_1/U134  ( .ZN(\MCD/adsel_1/n4356 ), .A(
        \stream3[45] ), .B(\MCD/adsel_1/n4355 ) );
    snl_nand02x1 \MCD/adsel_1/U108  ( .ZN(\MCD/adsel_1/n4339 ), .A(
        \MCD/adsel_1/n4337 ), .B(\MCD/adsel_1/n4340 ) );
    snl_invx05 \MCD/adsel_1/U141  ( .ZN(\MCD/adsel_1/n4322 ), .A(\stream3[48] 
        ) );
    snl_nand02x1 \MCD/adsel_1/U166  ( .ZN(\MCD/adsel_1/n4324 ), .A(
        \MCD/adsel_1/n4366 ), .B(\MCD/adsel_1/n4365 ) );
    snl_invx05 \MCD/adsel_1/U148  ( .ZN(\MCD/adsel_1/n4359 ), .A(
        \MCD/adsel_1/n4357 ) );
    snl_oai013x0 \MCD/adsel_1/U153  ( .ZN(\MCD/adsel_1/n4363 ), .A(
        \MCD/adsel_1/n4352 ), .B(\MCD/adsel_1/n4362 ), .C(\MCD/adsel_1/n4333 ), 
        .D(\stream3[33] ) );
    snl_ffqrnx1 \MCD/adsel_1/ciff_reg  ( .Q(\MCD/adsel_1/ciff ), .D(pk_ciffh), 
        .RN(n10733), .CP(SCLK) );
    snl_invx05 \MCD/adsel_1/U101  ( .ZN(\MCD/adsel_1/n4333 ), .A(\stream3[34] 
        ) );
    snl_nor02x1 \MCD/adsel_1/U106  ( .ZN(\MCD/adsel_1/n4337 ), .A(
        \MCD/adsel_1/n4328 ), .B(\stream3[59] ) );
    snl_nor02x1 \MCD/adsel_1/U121  ( .ZN(\MCD/adsel_1/n4319 ), .A(
        \MCD/adsel_1/n4345 ), .B(\MCD/adsel_1/n4288 ) );
    snl_oai222x0 \MCD/adsel_1/U126  ( .ZN(\MCD/adsel_1/n4348 ), .A(
        \MCD/adsel_1/bacc ), .B(\MCD/adsel_1/n4335 ), .C(\MCD/adsel_1/n4302 ), 
        .D(\MCD/adsel_1/n4336 ), .E(pk_sign_h), .F(\stream3[34] ) );
    snl_nand02x1 \MCD/adsel_1/U168  ( .ZN(\MCD/adsel_1/n4353 ), .A(ph_ioselh), 
        .B(\pk_stat_h[18] ) );
    snl_aoi113x0 \MCD/adsel_1/U91  ( .ZN(\MCD/adsel_1/n4326 ), .A(
        \stream3[41] ), .B(\MCD/adsel_1/n4323 ), .C(\MCD/adsel_1/n4327 ), .D(
        \MCD/adsel_1/n4320 ), .E(\MCD/adsel_1/n4314 ) );
    snl_nand13x1 \MCD/adsel_1/U98  ( .ZN(\MCD/adsel_1/n4287 ), .A(ph_saexe_sth
        ), .B(po_ptrsel_h), .C(ph_stage_ah) );
    snl_aoi022x1 \MCD/adsel_1/U128  ( .ZN(\MCD/adsel_1/n4350 ), .A(
        \MCD/adsel_1/n4303 ), .B(\stream3[32] ), .C(\MCD/adsel_1/bacc ), .D(
        \MCD/adsel_1/n4334 ) );
    snl_oai122x0 \MCD/adsel_1/U154  ( .ZN(\MCD/adsel_1/n4340 ), .A(
        \MCD/adsel_1/n4335 ), .B(\MCD/adsel_1/n4350 ), .C(\stream3[34] ), .D(
        \MCD/adsel_1/n4351 ), .E(\MCD/adsel_1/n4363 ) );
    snl_oai012x1 \MCD/adsel_1/U146  ( .ZN(\MCD/adsel_1/n4297 ), .A(
        \MCD/adsel_1/n4359 ), .B(\MCD/adsel_1/n4307 ), .C(ph_stage_ah) );
    snl_invx05 \MCD/adsel_1/U161  ( .ZN(\MCD/adsel_1/n4301 ), .A(po_sprtrs_h)
         );
    snl_and02x1 \MCD/adsel_1/U114  ( .Z(\MCD/adsel_1/n4305 ), .A(\stream3[41] 
        ), .B(\MCD/adsel_1/n4323 ) );
    snl_nor02x1 \MCD/adsel_1/U133  ( .ZN(\MCD/adsel_1/n4311 ), .A(
        \MCD/adsel_1/n4355 ), .B(\MCD/adsel_1/n4338 ) );
    snl_oai022x1 \MCD/adsel_1/U75  ( .ZN(po_dprtrs_h), .A(\MCD/adsel_1/n4291 ), 
        .B(\MCD/adsel_1/n4292 ), .C(\MCD/adsel_1/n4293 ), .D(
        \MCD/adsel_1/n4294 ) );
    snl_aoi012x1 \MCD/adsel_1/U82  ( .ZN(\MCD/adsel_1/n4304 ), .A(
        \stream3[32] ), .B(\MCD/adsel_1/n4303 ), .C(\stream3[33] ) );
    snl_invx05 \MCD/adsel_1/U99  ( .ZN(\MCD/adsel_1/n4288 ), .A(\stream3[40] )
         );
    snl_oai122x0 \MCD/adsel_1/U155  ( .ZN(\MCD/adsel_1/n4344 ), .A(
        \MCD/adsel_1/n4335 ), .B(\MCD/adsel_1/n4342 ), .C(\stream3[34] ), .D(
        \MCD/adsel_1/n4304 ), .E(\MCD/adsel_1/n4364 ) );
    snl_invx05 \MCD/adsel_1/U107  ( .ZN(\MCD/adsel_1/n4338 ), .A(\stream3[47] 
        ) );
    snl_aoi012x1 \MCD/adsel_1/U120  ( .ZN(\MCD/adsel_1/n4318 ), .A(stage_b), 
        .B(\MCD/adsel_1/n4299 ), .C(ph_exstgb_h) );
    snl_and02x1 \MCD/adsel_1/U115  ( .Z(\MCD/adsel_1/n4306 ), .A(\stream3[43] 
        ), .B(\MCD/adsel_1/n4310 ) );
    snl_aoi022x1 \MCD/adsel_1/U132  ( .ZN(\MCD/adsel_1/n4296 ), .A(
        \MCD/adsel_1/n4330 ), .B(\stream3[58] ), .C(\stream3[57] ), .D(
        \MCD/adsel_1/n4328 ) );
    snl_aoi223x0 \MCD/adsel_1/U90  ( .ZN(\MCD/adsel_1/n4284 ), .A(
        \MCD/adsel_1/n4321 ), .B(\MCD/adsel_1/n4322 ), .C(\MCD/adsel_1/n4323 ), 
        .D(po_mode01_h), .E(\MCD/adsel_1/n4324 ), .F(\MCD/adsel_1/n4310 ), .G(
        \MCD/adsel_1/n4325 ) );
    snl_invx05 \MCD/adsel_1/U97  ( .ZN(\MCD/adsel_1/n4299 ), .A(ph_stage_ah)
         );
    snl_nand03x0 \MCD/adsel_1/U109  ( .ZN(\MCD/adsel_1/n4308 ), .A(po_mode01_h
        ), .B(\MCD/adsel_1/n4338 ), .C(\stream3[46] ) );
    snl_aoi022x1 \MCD/adsel_1/U129  ( .ZN(\MCD/adsel_1/n4351 ), .A(
        \MCD/adsel_1/ciff ), .B(\stream3[32] ), .C(pk_sign_h), .D(
        \MCD/adsel_1/n4334 ) );
    snl_nand02x1 \MCD/adsel_1/U147  ( .ZN(\MCD/adsel_1/n4357 ), .A(
        \MCD/adsel_1/n4360 ), .B(\MCD/adsel_1/n4361 ) );
    snl_invx05 \MCD/adsel_1/U160  ( .ZN(\MCD/adsel_1/n4316 ), .A(
        \MCD/adsel_1/n4318 ) );
    snl_invx05 \MCD/adsel_1/U140  ( .ZN(\MCD/adsel_1/n4323 ), .A(
        \MCD/adsel_1/n4343 ) );
    snl_aoi022x1 \MCD/adsel_1/U167  ( .ZN(\MCD/adsel_1/n4364 ), .A(
        \MCD/adsel_1/n4349 ), .B(\stream3[32] ), .C(\MCD/adsel_1/n4348 ), .D(
        \MCD/adsel_1/n4334 ) );
    snl_aoi013x0 \MCD/adsel_1/U85  ( .ZN(\MCD/adsel_1/n4298 ), .A(
        \MCD/adsel_1/n4310 ), .B(\stream3[46] ), .C(\MCD/adsel_1/n4311 ), .D(
        \MCD/adsel_1/n4312 ) );
    snl_invx05 \MCD/adsel_1/U100  ( .ZN(\MCD/adsel_1/n4328 ), .A(\stream3[58] 
        ) );
    snl_invx05 \MCD/adsel_1/U112  ( .ZN(\MCD/adsel_1/n4309 ), .A(\stream3[44] 
        ) );
    snl_nand02x1 \MCD/adsel_1/U135  ( .ZN(\MCD/adsel_1/n4346 ), .A(
        \MCD/adsel_1/n4301 ), .B(\MCD/adsel_1/n4357 ) );
    snl_aoi122x0 \MCD/adsel_1/U127  ( .ZN(\MCD/adsel_1/n4349 ), .A(ph_ioselh), 
        .B(\pk_stat_h[18] ), .C(\MCD/adsel_1/bacc ), .D(\MCD/adsel_1/ciff ), 
        .E(\MCD/adsel_1/n4336 ) );
    snl_nand04x0 \MCD/adsel_1/U149  ( .ZN(\MCD/adsel_1/n4300 ), .A(
        \MCD/adsel_1/n4323 ), .B(\stream3[44] ), .C(\MCD/adsel_1/n4356 ), .D(
        \MCD/adsel_1/n4316 ) );
    snl_aoi013x0 \MCD/adsel_1/U137  ( .ZN(\MCD/adsel_1/n4327 ), .A(
        \MCD/adsel_1/n4336 ), .B(\MCD/adsel_1/n4333 ), .C(\stream3[32] ), .D(
        \stream3[40] ) );
    snl_invx05 \MCD/adsel_1/U152  ( .ZN(\MCD/adsel_1/n4362 ), .A(
        \MCD/adsel_1/n4342 ) );
    snl_nor02x1 \MCD/adsel_1/U71  ( .ZN(po_imdselh), .A(ph_saexe_sth), .B(
        \MCD/adsel_1/n4286 ) );
    snl_nor03x0 \MCD/adsel_1/U76  ( .ZN(po_bitsrc_h), .A(\stream3[52] ), .B(
        \stream3[53] ), .C(\stream3[54] ) );
    snl_oai112x0 \MCD/adsel_1/U77  ( .ZN(po_oprtrs_h), .A(\MCD/adsel_1/n4295 ), 
        .B(\MCD/adsel_1/n4296 ), .C(\MCD/adsel_1/n4297 ), .D(
        \MCD/adsel_1/n4289 ) );
    snl_oai012x1 \MCD/adsel_1/U79  ( .ZN(po_sprtrs_h), .A(\MCD/adsel_1/n4298 ), 
        .B(\MCD/adsel_1/n4299 ), .C(\MCD/adsel_1/n4300 ) );
    snl_nor02x1 \MCD/adsel_1/U95  ( .ZN(po_mode01_h), .A(\stream3[58] ), .B(
        \stream3[59] ) );
    snl_invx05 \MCD/adsel_1/U110  ( .ZN(\MCD/adsel_1/n4341 ), .A(\stream3[45] 
        ) );
    snl_oai033x0 \MCD/adsel_1/U159  ( .ZN(\MCD/adsel_1/n4360 ), .A(
        \MCD/adsel_1/n4343 ), .B(\stream3[44] ), .C(\MCD/adsel_1/n4341 ), .D(
        \MCD/adsel_1/n4339 ), .E(\stream3[46] ), .F(\MCD/adsel_1/n4338 ) );
    snl_oa023x1 \MCD/adsel_1/U119  ( .Z(\MCD/adsel_1/n4315 ), .A(
        \MCD/adsel_1/n4346 ), .B(\MCD/adsel_1/n4313 ), .C(\MCD/adsel_1/n4299 ), 
        .D(\MCD/adsel_1/n4317 ), .E(\MCD/adsel_1/n4347 ) );
    snl_invx05 \MCD/adsel_1/U142  ( .ZN(\MCD/adsel_1/n4292 ), .A(
        \MCD/adsel_1/n4319 ) );
    snl_nand14x0 \MCD/adsel_1/U165  ( .ZN(\MCD/adsel_1/n4366 ), .A(
        \stream3[46] ), .B(\MCD/adsel_1/n4338 ), .C(\MCD/adsel_1/n4341 ), .D(
        \MCD/adsel_1/n4309 ) );
    snl_nand02x1 \MCD/adsel_1/U80  ( .ZN(po_trsset_h), .A(\MCD/adsel_1/n4301 ), 
        .B(\MCD/adsel_1/n4290 ) );
    snl_aoi013x0 \MCD/adsel_1/U87  ( .ZN(\MCD/adsel_1/n4294 ), .A(ph_stage_ah), 
        .B(\MCD/adsel_1/n4297 ), .C(\MCD/adsel_1/n4315 ), .D(
        \MCD/adsel_1/n4316 ) );
    snl_invx05 \MCD/adsel_1/U150  ( .ZN(po_sprlth), .A(\MCD/adsel_1/n4300 ) );
    snl_invx05 \MCD/adsel_1/U102  ( .ZN(\MCD/adsel_1/n4334 ), .A(\stream3[32] 
        ) );
    snl_xor2x0 \MCD/adsel_1/U125  ( .Z(\MCD/adsel_1/n4331 ), .A(
        \MCD/adsel_1/bacc ), .B(\stream3[50] ) );
    snl_invx05 \MCD/adsel_1/U105  ( .ZN(\MCD/adsel_1/n4336 ), .A(\stream3[33] 
        ) );
    snl_and23x0 \MCD/adsel_1/U122  ( .Z(po_wrdsrc_h), .A(\stream3[54] ), .B(
        \stream3[53] ), .C(\stream3[52] ) );
    snl_nor04x0 \MCD/adsel_1/U89  ( .ZN(\MCD/adsel_1/n4285 ), .A(
        \MCD/adsel_1/n4319 ), .B(\MCD/adsel_1/n4320 ), .C(\MCD/adsel_1/n4306 ), 
        .D(\MCD/adsel_1/n4305 ) );
    snl_invx05 \MCD/adsel_1/U139  ( .ZN(\MCD/adsel_1/n4310 ), .A(
        \MCD/adsel_1/n4339 ) );
    snl_nand04x0 \MCD/adsel_1/U157  ( .ZN(\MCD/adsel_1/n4361 ), .A(
        \stream3[33] ), .B(\MCD/adsel_1/n4354 ), .C(\MCD/adsel_1/n4334 ), .D(
        \MCD/adsel_1/n4333 ) );
    snl_aoi013x0 \MCD/adsel_1/U92  ( .ZN(\MCD/adsel_1/n4286 ), .A(
        \MCD/adsel_1/n4328 ), .B(\MCD/adsel_1/n4329 ), .C(\stream3[59] ), .D(
        \stream3[54] ) );
    snl_invx05 \MCD/adsel_1/U145  ( .ZN(\MCD/adsel_1/n4347 ), .A(
        \MCD/adsel_1/n4320 ) );
    snl_invx05 \MCD/adsel_1/U162  ( .ZN(\MCD/adsel_1/n4290 ), .A(po_dprtrs_h)
         );
    snl_ao1b1b3x0 \MCD/adsel_1/U117  ( .Z(\MCD/adsel_1/n4317 ), .A(
        \MCD/adsel_1/n4309 ), .B(\stream3[45] ), .C(\MCD/adsel_1/n4308 ), .D(
        ph_stage_ah), .E(\MCD/adsel_1/n4312 ) );
    snl_nor02x1 \MCD/adsel_1/U81  ( .ZN(\MCD/adsel_1/n4302 ), .A(pk_pcon31_h), 
        .B(\MCD/adsel_1/n4303 ) );
    snl_aoi022x1 \MCD/adsel_1/U130  ( .ZN(\MCD/adsel_1/n4352 ), .A(
        \MCD/adsel_1/n4353 ), .B(\stream3[32] ), .C(\MCD/adsel_1/n4354 ), .D(
        \MCD/adsel_1/n4334 ) );
    snl_invx05 \MCD/adsel_1/U138  ( .ZN(\MCD/adsel_1/n4358 ), .A(pk_pcon31_h)
         );
    snl_nand02x1 \MCD/adsel_1/U156  ( .ZN(\MCD/adsel_1/n4354 ), .A(
        \MCD/adsel_1/ciff ), .B(\MCD/adsel_1/n4358 ) );
    snl_nand02x1 \MCD/adsel_1/U104  ( .ZN(\MCD/adsel_1/n4335 ), .A(
        \stream3[34] ), .B(\MCD/adsel_1/n4336 ) );
    snl_nand14x0 \MCD/adsel_1/U116  ( .ZN(\MCD/adsel_1/n4345 ), .A(
        \stream3[43] ), .B(\stream3[41] ), .C(po_mode01_h), .D(
        \MCD/adsel_1/n4332 ) );
    snl_invx05 \MCD/adsel_1/U123  ( .ZN(\MCD/adsel_1/n4295 ), .A(\stream3[59] 
        ) );
    snl_ffqrnx1 \MCD/adsel_1/bacc_reg  ( .Q(\MCD/adsel_1/bacc ), .D(pk_bacch), 
        .RN(n10733), .CP(SCLK) );
    snl_and02x1 \MCD/adsel_1/U88  ( .Z(\MCD/adsel_1/n4291 ), .A(
        \MCD/adsel_1/n4317 ), .B(\MCD/adsel_1/n4318 ) );
    snl_aoi012x1 \MCD/adsel_1/U93  ( .ZN(\MCD/adsel_1/n4330 ), .A(
        \stream3[51] ), .B(\MCD/adsel_1/n4331 ), .C(\stream3[57] ) );
    snl_invx05 \MCD/adsel_1/U131  ( .ZN(\MCD/adsel_1/n4329 ), .A(\stream3[57] 
        ) );
    snl_invx05 \MCD/adsel_1/U94  ( .ZN(\MCD/adsel_1/n4332 ), .A(\stream3[42] )
         );
    snl_nor03x0 \MCD/adsel_1/U143  ( .ZN(\MCD/adsel_1/n4312 ), .A(
        \MCD/adsel_1/n4308 ), .B(\stream3[44] ), .C(\MCD/adsel_1/n4341 ) );
    snl_invx05 \MCD/adsel_1/U144  ( .ZN(\MCD/adsel_1/n4321 ), .A(\stream3[49] 
        ) );
    snl_oai023x0 \MCD/adsel_1/U163  ( .ZN(\MCD/adsel_1/n4325 ), .A(
        \MCD/adsel_1/n4355 ), .B(\stream3[46] ), .C(\stream3[47] ), .D(
        \stream3[51] ), .E(\stream3[50] ) );
    snl_invx05 \MCD/adsel_1/U158  ( .ZN(\MCD/adsel_1/n4355 ), .A(
        \MCD/adsel_1/n4361 ) );
    snl_or04x1 \MCD/adsel_1/U164  ( .Z(\MCD/adsel_1/n4365 ), .A(\stream3[49] ), 
        .B(\stream3[48] ), .C(\stream3[50] ), .D(\stream3[51] ) );
    snl_nand03x0 \MCD/adsel_1/U136  ( .ZN(\MCD/adsel_1/n4283 ), .A(po_wrdsrc_h
        ), .B(ph_stage_ah), .C(\stream3[55] ) );
    snl_and23x0 \MCD/adsel_1/U78  ( .Z(po_lwdsrc_h), .A(\stream3[54] ), .B(
        \stream3[52] ), .C(\stream3[53] ) );
    snl_aoi012x1 \MCD/adsel_1/U86  ( .ZN(\MCD/adsel_1/n4313 ), .A(
        \MCD/adsel_1/n4305 ), .B(\MCD/adsel_1/n4288 ), .C(\MCD/adsel_1/n4314 )
         );
    snl_invx05 \MCD/adsel_1/U103  ( .ZN(\MCD/adsel_1/n4303 ), .A(
        \MCD/adsel_1/ciff ) );
    snl_nand03x0 \MCD/adsel_1/U111  ( .ZN(\MCD/adsel_1/n4342 ), .A(
        \MCD/adsel_1/ciff ), .B(\stream3[32] ), .C(\MCD/adsel_1/bacc ) );
    snl_oa012x1 \MCD/adsel_1/U124  ( .Z(\MCD/adsel_1/n4289 ), .A(
        \MCD/adsel_1/n4318 ), .B(\MCD/adsel_1/n4326 ), .C(\MCD/adsel_1/n4315 )
         );
    snl_nor02x1 \MCD/adsel_1/U118  ( .ZN(\MCD/adsel_1/n4320 ), .A(
        \MCD/adsel_1/n4345 ), .B(\stream3[40] ) );
    snl_and02x1 \MCD/adsel_1/U151  ( .Z(\MCD/adsel_1/n4314 ), .A(
        \MCD/adsel_1/n4306 ), .B(\MCD/adsel_1/n4332 ) );
    snl_oai022x1 \LBUS/phsdlt_1/U25  ( .ZN(\LBUS/phsdlt_1/nrt[2] ), .A(
        \LBUS/srdalth ), .B(\LBUS/phsdlt_1/n1012 ), .C(\LBUS/phsdlt_1/n1013 ), 
        .D(\LBUS/phsdlt_1/n1014 ) );
    snl_aoi012x1 \LBUS/phsdlt_1/U26  ( .ZN(\LBUS/phsdlt_1/nrt[1] ), .A(
        \LBUS/phsdlt_1/n1012 ), .B(\LBUS/phsdlt_1/n1015 ), .C(\LBUS/srdalth )
         );
    snl_invx05 \LBUS/phsdlt_1/U28  ( .ZN(\LBUS/phsdlt_1/n1013 ), .A(ph_bit_h)
         );
    snl_oai022x1 \LBUS/phsdlt_1/U27  ( .ZN(\LBUS/phsdlt_1/nrt[0] ), .A(
        \LBUS/srdalth ), .B(\LBUS/phsdlt_1/n1015 ), .C(ph_bit_h), .D(
        \LBUS/phsdlt_1/n1014 ) );
    snl_ffqrnx1 \LBUS/phsdlt_1/irt_reg[1]  ( .Q(\LBUS/srdalth ), .D(
        \LBUS/phsdlt_1/nrt[1] ), .RN(n10734), .CP(SCLK) );
    snl_nand03x0 \LBUS/phsdlt_1/U29  ( .ZN(\LBUS/phsdlt_1/n1014 ), .A(
        \LBUS/phsdlt_1/n1015 ), .B(\LBUS/phsdlt_1/n1012 ), .C(ph_lpdilth) );
    snl_invx05 \LBUS/phsdlt_1/U30  ( .ZN(\LBUS/phsdlt_1/n1012 ), .A(
        ph_btsrdaselh) );
    snl_ffqrnx1 \LBUS/phsdlt_1/irt_reg[0]  ( .Q(ph_wdsrdaselh), .D(
        \LBUS/phsdlt_1/nrt[0] ), .RN(n10734), .CP(SCLK) );
    snl_ffqrnx1 \LBUS/phsdlt_1/irt_reg[2]  ( .Q(ph_btsrdaselh), .D(
        \LBUS/phsdlt_1/nrt[2] ), .RN(n10734), .CP(SCLK) );
    snl_invx05 \LBUS/phsdlt_1/U31  ( .ZN(\LBUS/phsdlt_1/n1015 ), .A(
        ph_wdsrdaselh) );
    snl_bufx1 \CONS/phsegsel_1/U21  ( .Z(\CONS/phsegsel_1/n328 ), .A(
        ph_tprsel_h) );
    snl_and24x0 \CONS/phsegsel_1/U22  ( .Z(ph_ioselh), .A(\stream3[30] ), .B(
        \stream3[29] ), .C(\stream3[31] ), .D(\stream3[28] ) );
    snl_aoi222x0 \CONS/phsegsel_1/U26  ( .ZN(\CONS/phsegsel_1/n336 ), .A(
        ph_srcadr1_h), .B(\pk_sra1_h[31] ), .C(\CONS/phsegsel_1/n328 ), .D(
        \pk_trba_h[31] ), .E(ph_srcadr2_h), .F(\pk_sra2_h[31] ) );
    snl_aoi222x0 \CONS/phsegsel_1/U28  ( .ZN(\CONS/phsegsel_1/n333 ), .A(
        \pk_sra1_h[30] ), .B(ph_srcadr1_h), .C(\pk_trba_h[30] ), .D(
        \CONS/phsegsel_1/n328 ), .E(\pk_sra2_h[30] ), .F(ph_srcadr2_h) );
    snl_aoi222x0 \CONS/phsegsel_1/U33  ( .ZN(\CONS/phsegsel_1/n334 ), .A(
        \stream3[28] ), .B(ph_oprtrs_h), .C(\pk_spr_h[28] ), .D(ph_sprtrs_h), 
        .E(\pk_dpr_h[28] ), .F(ph_dprtrs_h) );
    snl_and02x1 \CONS/phsegsel_1/U34  ( .Z(ph_obmselh), .A(
        \CONS/phsegsel_1/n337 ), .B(\CONS/phsegsel_1/n336 ) );
    snl_aoi222x0 \CONS/phsegsel_1/U27  ( .ZN(\CONS/phsegsel_1/n337 ), .A(
        ph_oprtrs_h), .B(\stream3[31] ), .C(ph_sprtrs_h), .D(\pk_spr_h[31] ), 
        .E(ph_dprtrs_h), .F(\pk_dpr_h[31] ) );
    snl_aoi222x0 \CONS/phsegsel_1/U29  ( .ZN(\CONS/phsegsel_1/n332 ), .A(
        \stream3[30] ), .B(ph_oprtrs_h), .C(\pk_spr_h[30] ), .D(ph_sprtrs_h), 
        .E(\pk_dpr_h[30] ), .F(ph_dprtrs_h) );
    snl_aoi222x0 \CONS/phsegsel_1/U32  ( .ZN(\CONS/phsegsel_1/n335 ), .A(
        \pk_sra1_h[28] ), .B(ph_srcadr1_h), .C(\pk_trba_h[28] ), .D(
        \CONS/phsegsel_1/n328 ), .E(\pk_sra2_h[28] ), .F(ph_srcadr2_h) );
    snl_nor02x1 \CONS/phsegsel_1/U23  ( .ZN(ph_mmbselh), .A(ph_obmselh), .B(
        \CONS/phsegsel_1/n329 ) );
    snl_and12x1 \CONS/phsegsel_1/U24  ( .Z(ph_extselh), .A(ph_obmselh), .B(
        \CONS/phsegsel_1/n329 ) );
    snl_aoi222x0 \CONS/phsegsel_1/U25  ( .ZN(\CONS/phsegsel_1/n329 ), .A(
        \CONS/phsegsel_1/n330 ), .B(\CONS/phsegsel_1/n331 ), .C(
        \CONS/phsegsel_1/n332 ), .D(\CONS/phsegsel_1/n333 ), .E(
        \CONS/phsegsel_1/n334 ), .F(\CONS/phsegsel_1/n335 ) );
    snl_aoi222x0 \CONS/phsegsel_1/U30  ( .ZN(\CONS/phsegsel_1/n331 ), .A(
        \pk_sra1_h[29] ), .B(ph_srcadr1_h), .C(\pk_trba_h[29] ), .D(
        \CONS/phsegsel_1/n328 ), .E(\pk_sra2_h[29] ), .F(ph_srcadr2_h) );
    snl_aoi222x0 \CONS/phsegsel_1/U31  ( .ZN(\CONS/phsegsel_1/n330 ), .A(
        \stream3[29] ), .B(ph_oprtrs_h), .C(\pk_spr_h[29] ), .D(ph_sprtrs_h), 
        .E(\pk_dpr_h[29] ), .F(ph_dprtrs_h) );
    snl_mux21x1 \ADOSEL/seladr_1/U10  ( .Z(LOUT[7]), .A(\pgsadrh[7] ), .B(
        \pgmuxout[7] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U12  ( .Z(LOUT[5]), .A(\pgsadrh[5] ), .B(
        \pgmuxout[5] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U13  ( .Z(LOUT[4]), .A(\pgsadrh[4] ), .B(
        \pgmuxout[4] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U14  ( .Z(LOUT[3]), .A(\pgsadrh[3] ), .B(
        \pgmuxout[3] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U15  ( .Z(LOUT[2]), .A(\pgsadrh[2] ), .B(
        \pgmuxout[2] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U17  ( .Z(LOUT[0]), .A(\pgsadrh[0] ), .B(
        \pgmuxout[0] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U11  ( .Z(LOUT[6]), .A(\pgsadrh[6] ), .B(
        \pgmuxout[6] ), .S(ph_ldaoutenh1) );
    snl_mux21x1 \ADOSEL/seladr_1/U16  ( .Z(LOUT[1]), .A(\pgsadrh[1] ), .B(
        \pgmuxout[1] ), .S(ph_ldaoutenh1) );
    snl_and02x1 \LBUS/ldoecnt_1/U8  ( .Z(ph_ldaoutenh1), .A(ph_lbwrh), .B(
        \LBUS/temp[3] ) );
    snl_ao022x1 \REG_2/SATIME/U33  ( .Z(\REG_2/SATIME/count97[20] ), .A(
        \pk_stdat[20] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[20] ), .D(\REG_2/SATIME/n228 ) );
    snl_nor02x1 \REG_2/SATIME/U54  ( .ZN(\REG_2/SATIME/ph_timouth117 ), .A(
        \REG_2/SATIME/count[19] ), .B(\REG_2/SATIME/n229 ) );
    snl_invx05 \REG_2/SATIME/U73  ( .ZN(\REG_2/SATIME/n246 ), .A(
        \REG_2/SATIME/count[8] ) );
    snl_invx05 \REG_2/SATIME/U68  ( .ZN(\REG_2/SATIME/n232 ), .A(
        \REG_2/SATIME/count[1] ) );
    snl_oai112x0 \REG_2/SATIME/U96  ( .ZN(\REG_2/SATIME/n249 ), .A(
        \REG_2/SATIME/n230 ), .B(\REG_2/SATIME/n235 ), .C(\REG_2/SATIME/n257 ), 
        .D(\REG_2/SATIME/count[9] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[6]  ( .Q(\REG_2/SATIME/count[6] ), .D(
        \REG_2/SATIME/count97[6] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/dda1_reg  ( .Q(\REG_2/SATIME/dda1 ), .D(
        \pk_sati_h[1] ), .CP(SCLK) );
    snl_ao022x1 \REG_2/SATIME/U34  ( .Z(\REG_2/SATIME/count97[19] ), .A(
        \pk_stdat[19] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[19] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U41  ( .Z(\REG_2/SATIME/count97[12] ), .A(
        \pk_stdat[12] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[12] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U46  ( .Z(\REG_2/SATIME/count97[7] ), .A(
        \pk_stdat[7] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[7] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_and08x1 \REG_2/SATIME/U61  ( .Z(\REG_2/SATIME/n252 ), .A(
        \REG_2/SATIME/n253 ), .B(\REG_2/SATIME/n254 ), .C(\REG_2/SATIME/n251 ), 
        .D(\REG_2/SATIME/n244 ), .E(\REG_2/SATIME/n255 ), .F(
        \REG_2/SATIME/n256 ), .G(\REG_2/SATIME/n257 ), .H(\REG_2/SATIME/n258 )
         );
    snl_aoi022x1 \REG_2/SATIME/U84  ( .ZN(\REG_2/SATIME/n261 ), .A(
        \REG_2/SATIME/n242 ), .B(\REG_2/SATIME/count[0] ), .C(
        \REG_2/SATIME/n248 ), .D(\REG_2/SATIME/n254 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[2]  ( .Q(\REG_2/SATIME/count[2] ), .D(
        \REG_2/SATIME/count97[2] ), .CP(SCLK) );
    snl_invx05 \REG_2/SATIME/U101  ( .ZN(\REG_2/SATIME/n245 ), .A(
        \REG_2/SATIME/n236 ) );
    snl_nand13x1 \REG_2/SATIME/U66  ( .ZN(\REG_2/SATIME/n233 ), .A(
        \REG_2/SATIME/count[17] ), .B(\REG_2/SATIME/count[7] ), .C(
        \REG_2/SATIME/count[3] ) );
    snl_aoi022x1 \REG_2/SATIME/U83  ( .ZN(\REG_2/SATIME/n237 ), .A(
        \REG_2/SATIME/n238 ), .B(\REG_2/SATIME/count[6] ), .C(
        \REG_2/SATIME/n241 ), .D(\REG_2/SATIME/n255 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[0]  ( .Q(\REG_2/SATIME/count[0] ), .D(
        \REG_2/SATIME/count97[0] ), .CP(SCLK) );
    snl_nand03x0 \REG_2/SATIME/U98  ( .ZN(\REG_2/SATIME/n260 ), .A(
        \REG_2/SATIME/count[14] ), .B(\REG_2/SATIME/n266 ), .C(
        \REG_2/SATIME/count[13] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[9]  ( .Q(\REG_2/SATIME/count[9] ), .D(
        \REG_2/SATIME/count97[9] ), .CP(SCLK) );
    snl_ao022x1 \REG_2/SATIME/U35  ( .Z(\REG_2/SATIME/count97[18] ), .A(
        \pk_stdat[18] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[18] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U48  ( .Z(\REG_2/SATIME/count97[5] ), .A(
        \pk_stdat[5] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[5] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[4]  ( .Q(\REG_2/SATIME/count[4] ), .D(
        \REG_2/SATIME/count97[4] ), .CP(SCLK) );
    snl_ao022x1 \REG_2/SATIME/U53  ( .Z(\REG_2/SATIME/count97[0] ), .A(
        \pk_stdat[0] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[0] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_muxi21x1 \REG_2/SATIME/U91  ( .ZN(\REG_2/SATIME/n229 ), .A(
        \REG_2/SATIME/n252 ), .B(\REG_2/SATIME/n259 ), .S(
        \REG_2/SATIME/count[12] ) );
    snl_invx05 \REG_2/SATIME/U74  ( .ZN(\REG_2/SATIME/n251 ), .A(
        \REG_2/SATIME/count[5] ) );
    snl_invx05 \REG_2/SATIME/U99  ( .ZN(\REG_2/SATIME/n254 ), .A(
        \REG_2/SATIME/count[0] ) );
    snl_ao022x1 \REG_2/SATIME/U36  ( .Z(\REG_2/SATIME/count97[17] ), .A(
        \pk_stdat[17] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[17] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U37  ( .Z(\REG_2/SATIME/count97[16] ), .A(
        \pk_stdat[16] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[16] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U39  ( .Z(\REG_2/SATIME/count97[14] ), .A(
        \pk_stdat[14] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[14] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U40  ( .Z(\REG_2/SATIME/count97[13] ), .A(
        \pk_stdat[13] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[13] ), .D(\REG_2/SATIME/n228 ) );
    snl_and02x1 \REG_2/SATIME/U82  ( .Z(\REG_2/SATIME/n227 ), .A(
        \pk_rwrit_h[1] ), .B(\REG_2/SATIME/n267 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[18]  ( .Q(\REG_2/SATIME/count[18] ), .D(
        \REG_2/SATIME/count97[18] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/count_reg[11]  ( .Q(\REG_2/SATIME/count[11] ), .D(
        \REG_2/SATIME/count97[11] ), .CP(SCLK) );
    snl_ao022x1 \REG_2/SATIME/U47  ( .Z(\REG_2/SATIME/count97[6] ), .A(
        \pk_stdat[6] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[6] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U49  ( .Z(\REG_2/SATIME/count97[4] ), .A(
        \pk_stdat[4] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[4] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U52  ( .Z(\REG_2/SATIME/count97[1] ), .A(
        \pk_stdat[1] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[1] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_nand04x0 \REG_2/SATIME/U67  ( .ZN(\REG_2/SATIME/n234 ), .A(
        \REG_2/SATIME/dda1 ), .B(\REG_2/SATIME/count[2] ), .C(
        \REG_2/SATIME/count[6] ), .D(\REG_2/SATIME/n263 ) );
    snl_invx05 \REG_2/SATIME/U75  ( .ZN(\REG_2/SATIME/n250 ), .A(
        \REG_2/SATIME/count[4] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[15]  ( .Q(\REG_2/SATIME/count[15] ), .D(
        \REG_2/SATIME/count97[15] ), .CP(SCLK) );
    snl_nand04x0 \REG_2/SATIME/U90  ( .ZN(\REG_2/SATIME/n276 ), .A(
        \REG_2/SATIME/n264 ), .B(\REG_2/SATIME/count[10] ), .C(
        \REG_2/SATIME/count[20] ), .D(\REG_2/SATIME/n277 ) );
    snl_nor04x0 \REG_2/SATIME/U55  ( .ZN(\REG_2/SATIME/n230 ), .A(
        \REG_2/SATIME/n231 ), .B(\REG_2/SATIME/n232 ), .C(\REG_2/SATIME/n233 ), 
        .D(\REG_2/SATIME/n234 ) );
    snl_invx05 \REG_2/SATIME/U69  ( .ZN(\REG_2/SATIME/n263 ), .A(
        \REG_2/SATIME/dda0 ) );
    snl_invx05 \REG_2/SATIME/U72  ( .ZN(\REG_2/SATIME/n244 ), .A(
        \REG_2/SATIME/count[9] ) );
    snl_nor03x0 \REG_2/SATIME/U97  ( .ZN(\REG_2/SATIME/n247 ), .A(
        \REG_2/SATIME/count[5] ), .B(\REG_2/SATIME/count[3] ), .C(
        \REG_2/SATIME/count[4] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[17]  ( .Q(\REG_2/SATIME/count[17] ), .D(
        \REG_2/SATIME/count97[17] ), .CP(SCLK) );
    snl_nor04x0 \REG_2/SATIME/U60  ( .ZN(\REG_2/SATIME/n248 ), .A(
        \REG_2/SATIME/n249 ), .B(\REG_2/SATIME/n250 ), .C(\REG_2/SATIME/n246 ), 
        .D(\REG_2/SATIME/n251 ) );
    snl_invx05 \REG_2/SATIME/U100  ( .ZN(\REG_2/SATIME/n243 ), .A(
        \REG_2/SATIME/n234 ) );
    snl_and03x1 \REG_2/SATIME/U57  ( .Z(\REG_2/SATIME/n238 ), .A(
        \REG_2/SATIME/count[17] ), .B(\REG_2/SATIME/n239 ), .C(
        \REG_2/SATIME/n240 ) );
    snl_nand03x0 \REG_2/SATIME/U85  ( .ZN(\REG_2/SATIME/n269 ), .A(
        \REG_2/SATIME/count[4] ), .B(\REG_2/SATIME/n240 ), .C(
        \REG_2/SATIME/count[14] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[20]  ( .Q(\REG_2/SATIME/count[20] ), .D(
        \REG_2/SATIME/count97[20] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/count_reg[13]  ( .Q(\REG_2/SATIME/count[13] ), .D(
        \REG_2/SATIME/count97[13] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/dda2_reg  ( .Q(\REG_2/SATIME/dda2 ), .D(
        \pk_sati_h[2] ), .CP(SCLK) );
    snl_nor02x1 \REG_2/SATIME/U70  ( .ZN(\REG_2/SATIME/n240 ), .A(
        \REG_2/SATIME/n263 ), .B(\REG_2/SATIME/count[3] ) );
    snl_ao022x1 \REG_2/SATIME/U42  ( .Z(\REG_2/SATIME/count97[11] ), .A(
        \pk_stdat[11] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[11] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U45  ( .Z(\REG_2/SATIME/count97[8] ), .A(
        \pk_stdat[8] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[8] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_invx05 \REG_2/SATIME/U79  ( .ZN(\REG_2/SATIME/n266 ), .A(
        \REG_2/SATIME/count[20] ) );
    snl_or03x1 \REG_2/SATIME/U95  ( .Z(\REG_2/SATIME/n231 ), .A(
        \REG_2/SATIME/count[15] ), .B(\REG_2/SATIME/count[16] ), .C(
        \REG_2/SATIME/dda2 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[12]  ( .Q(\REG_2/SATIME/count[12] ), .D(
        \REG_2/SATIME/count97[12] ), .CP(SCLK) );
    snl_nand03x0 \REG_2/SATIME/U87  ( .ZN(\REG_2/SATIME/n271 ), .A(
        \REG_2/SATIME/count[1] ), .B(\REG_2/SATIME/n250 ), .C(
        \REG_2/SATIME/n264 ) );
    snl_and34x0 \REG_2/SATIME/U62  ( .Z(\REG_2/SATIME/n259 ), .A(
        \REG_2/SATIME/n260 ), .B(\REG_2/SATIME/n261 ), .C(\REG_2/SATIME/n262 ), 
        .D(\REG_2/SATIME/count[11] ) );
    snl_invx05 \REG_2/SATIME/U65  ( .ZN(\REG_2/SATIME/n239 ), .A(
        \REG_2/SATIME/count[7] ) );
    snl_muxi21x1 \REG_2/SATIME/U102  ( .ZN(\REG_2/SATIME/n273 ), .A(
        \REG_2/SATIME/n269 ), .B(\REG_2/SATIME/n270 ), .S(
        \REG_2/SATIME/count[13] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[16]  ( .Q(\REG_2/SATIME/count[16] ), .D(
        \REG_2/SATIME/count97[16] ), .CP(SCLK) );
    snl_invx05 \REG_2/SATIME/U105  ( .ZN(\REG_2/SATIME/n268 ), .A(\REG_2/n435 
        ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[14]  ( .Q(\REG_2/SATIME/count[14] ), .D(
        \REG_2/SATIME/count97[14] ), .CP(SCLK) );
    snl_nor02x1 \REG_2/SATIME/U80  ( .ZN(\REG_2/SATIME/n267 ), .A(ph_timouth), 
        .B(\REG_2/SATIME/n268 ) );
    snl_ao022x1 \REG_2/SATIME/U50  ( .Z(\REG_2/SATIME/count97[3] ), .A(
        \pk_stdat[3] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[3] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_and08x1 \REG_2/SATIME/U59  ( .Z(\REG_2/SATIME/n242 ), .A(
        \REG_2/SATIME/n243 ), .B(\REG_2/SATIME/n244 ), .C(
        \REG_2/SATIME/count[17] ), .D(\REG_2/SATIME/count[18] ), .E(
        \REG_2/SATIME/n245 ), .F(\REG_2/SATIME/n246 ), .G(\REG_2/SATIME/n239 ), 
        .H(\REG_2/SATIME/n247 ) );
    snl_invx05 \REG_2/SATIME/U77  ( .ZN(\REG_2/SATIME/n262 ), .A(
        \REG_2/SATIME/count[10] ) );
    snl_nand04x0 \REG_2/SATIME/U89  ( .ZN(\REG_2/SATIME/n274 ), .A(
        \REG_2/SATIME/n275 ), .B(\REG_2/SATIME/n266 ), .C(\REG_2/SATIME/n262 ), 
        .D(\REG_2/SATIME/n246 ) );
    snl_nor02x1 \REG_2/SATIME/U92  ( .ZN(\REG_2/SATIME/n265 ), .A(
        \REG_2/SATIME/count[13] ), .B(\REG_2/SATIME/count[14] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[10]  ( .Q(\REG_2/SATIME/count[10] ), .D(
        \REG_2/SATIME/count97[10] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/count_reg[19]  ( .Q(\REG_2/SATIME/count[19] ), .D(
        \REG_2/SATIME/count97[19] ), .CP(SCLK) );
    snl_nor02x1 \REG_2/SATIME/U58  ( .ZN(\REG_2/SATIME/n241 ), .A(
        \REG_2/SATIME/dda0 ), .B(\REG_2/SATIME/n233 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[5]  ( .Q(\REG_2/SATIME/count[5] ), .D(
        \REG_2/SATIME/count97[5] ), .CP(SCLK) );
    snl_ao022x1 \REG_2/SATIME/U38  ( .Z(\REG_2/SATIME/count97[15] ), .A(
        \pk_stdat[15] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[15] ), .D(\REG_2/SATIME/n228 ) );
    snl_ao022x1 \REG_2/SATIME/U43  ( .Z(\REG_2/SATIME/count97[10] ), .A(
        \pk_stdat[10] ), .B(\REG_2/SATIME/n227 ), .C(
        \REG_2/SATIME/count145[10] ), .D(\REG_2/SATIME/n228 ) );
    snl_invx05 \REG_2/SATIME/U64  ( .ZN(\REG_2/SATIME/n253 ), .A(
        \REG_2/SATIME/count[2] ) );
    snl_and13x1 \REG_2/SATIME/U81  ( .Z(\REG_2/SATIME/n228 ), .A(
        \pk_rwrit_h[1] ), .B(\REG_2/SATIME/n267 ), .C(ph_timsth) );
    snl_muxi21x1 \REG_2/SATIME/U104  ( .ZN(\REG_2/SATIME/n256 ), .A(
        \REG_2/SATIME/n274 ), .B(\REG_2/SATIME/n276 ), .S(\REG_2/SATIME/dda2 )
         );
    snl_ao022x1 \REG_2/SATIME/U51  ( .Z(\REG_2/SATIME/count97[2] ), .A(
        \pk_stdat[2] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[2] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_invx05 \REG_2/SATIME/U76  ( .ZN(\REG_2/SATIME/n257 ), .A(
        \REG_2/SATIME/count[18] ) );
    snl_nand14x0 \REG_2/SATIME/U88  ( .ZN(\REG_2/SATIME/n272 ), .A(
        \REG_2/SATIME/dda1 ), .B(\REG_2/SATIME/n273 ), .C(\REG_2/SATIME/n239 ), 
        .D(\REG_2/SATIME/n232 ) );
    snl_nor04x0 \REG_2/SATIME/U93  ( .ZN(\REG_2/SATIME/n277 ), .A(
        \REG_2/SATIME/count[1] ), .B(\REG_2/SATIME/count[16] ), .C(
        \REG_2/SATIME/n246 ), .D(\REG_2/SATIME/n250 ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[1]  ( .Q(\REG_2/SATIME/count[1] ), .D(
        \REG_2/SATIME/count97[1] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/dda0_reg  ( .Q(\REG_2/SATIME/dda0 ), .D(
        \pk_sati_h[0] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/count_reg[8]  ( .Q(\REG_2/SATIME/count[8] ), .D(
        \REG_2/SATIME/count97[8] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/count_reg[3]  ( .Q(\REG_2/SATIME/count[3] ), .D(
        \REG_2/SATIME/count97[3] ), .CP(SCLK) );
    snl_ffqx1 \REG_2/SATIME/ph_timouth_reg  ( .Q(ph_timouth), .D(
        \REG_2/SATIME/ph_timouth117 ), .CP(SCLK) );
    snl_ao022x1 \REG_2/SATIME/U44  ( .Z(\REG_2/SATIME/count97[9] ), .A(
        \pk_stdat[9] ), .B(\REG_2/SATIME/n227 ), .C(\REG_2/SATIME/count145[9] 
        ), .D(\REG_2/SATIME/n228 ) );
    snl_nor04x0 \REG_2/SATIME/U56  ( .ZN(\REG_2/SATIME/n235 ), .A(
        \REG_2/SATIME/dda1 ), .B(\REG_2/SATIME/count[2] ), .C(
        \REG_2/SATIME/n236 ), .D(\REG_2/SATIME/n237 ) );
    snl_nor03x0 \REG_2/SATIME/U94  ( .ZN(\REG_2/SATIME/n258 ), .A(
        \REG_2/SATIME/count[17] ), .B(\REG_2/SATIME/count[11] ), .C(
        \REG_2/SATIME/count[15] ) );
    snl_nand04x0 \REG_2/SATIME/U71  ( .ZN(\REG_2/SATIME/n236 ), .A(
        \REG_2/SATIME/dda2 ), .B(\REG_2/SATIME/count[16] ), .C(
        \REG_2/SATIME/count[15] ), .D(\REG_2/SATIME/n232 ) );
    snl_invx05 \REG_2/SATIME/U63  ( .ZN(\REG_2/SATIME/n255 ), .A(
        \REG_2/SATIME/count[6] ) );
    snl_and04x1 \REG_2/SATIME/U78  ( .Z(\REG_2/SATIME/n264 ), .A(
        \REG_2/SATIME/n240 ), .B(\REG_2/SATIME/count[7] ), .C(
        \REG_2/SATIME/n265 ), .D(\REG_2/SATIME/dda1 ) );
    snl_nand14x0 \REG_2/SATIME/U86  ( .ZN(\REG_2/SATIME/n270 ), .A(
        \REG_2/SATIME/count[14] ), .B(\REG_2/SATIME/count[3] ), .C(
        \REG_2/SATIME/n250 ), .D(\REG_2/SATIME/n263 ) );
    snl_muxi21x1 \REG_2/SATIME/U103  ( .ZN(\REG_2/SATIME/n275 ), .A(
        \REG_2/SATIME/n272 ), .B(\REG_2/SATIME/n271 ), .S(
        \REG_2/SATIME/count[16] ) );
    snl_ffqx1 \REG_2/SATIME/count_reg[7]  ( .Q(\REG_2/SATIME/count[7] ), .D(
        \REG_2/SATIME/count97[7] ), .CP(SCLK) );
    snl_invx1 \SAEXE/RFIO/U224  ( .ZN(\SAEXE/RFIO/n386 ), .A(
        \SAEXE/RFIO/cnt4out[3] ) );
    snl_oai122x0 \SAEXE/RFIO/U231  ( .ZN(\SAEXE/RFIO/nfst[3] ), .A(
        \SAEXE/RFIO/n363 ), .B(\SAEXE/RFIO/n364 ), .C(\SAEXE/RFIO/n365 ), .D(
        \SAEXE/RFIO/n366 ), .E(\SAEXE/RFIO/n367 ) );
    snl_nor02x1 \SAEXE/RFIO/U238  ( .ZN(\SAEXE/RFIO/*cell*3735/U61/Z_0 ), .A(
        pgadrovfh), .B(\SAEXE/RFIO/n379 ) );
    snl_invx05 \SAEXE/RFIO/U256  ( .ZN(\SAEXE/RFIO/n377 ), .A(
        \SAEXE/RFIO/fst[2] ) );
    snl_invx05 \SAEXE/RFIO/U271  ( .ZN(\SAEXE/RFIO/n368 ), .A(
        \SAEXE/RFIO/cnt4out[2] ) );
    snl_invx05 \SAEXE/RFIO/U294  ( .ZN(\SAEXE/RFIO/n360 ), .A(
        \SAEXE/RFIO/n387 ) );
    snl_invx05 \SAEXE/RFIO/U304  ( .ZN(\SAEXE/RFIO/n404 ), .A(\pk_psae_h[7] )
         );
    snl_aoi223x0 \SAEXE/RFIO/U244  ( .ZN(\SAEXE/RFIO/n380 ), .A(
        \SAEXE/RFIO/n387 ), .B(\SAEXE/RFIO/n388 ), .C(\SAEXE/RFIO/cnt4out[3] ), 
        .D(\SAEXE/RFIO/n373 ), .E(\SAEXE/RFIO/n376 ), .F(\SAEXE/RFIO/n389 ), 
        .G(\SAEXE/RFIO/n390 ) );
    snl_and34x0 \SAEXE/RFIO/U286  ( .Z(\SAEXE/RFIO/rfin2h ), .A(\pk_psae_h[6] 
        ), .B(\SAEXE/RFIO/n404 ), .C(\pk_psae_h[5] ), .D(\pk_psae_h[4] ) );
    snl_invx05 \SAEXE/RFIO/U263  ( .ZN(\SAEXE/RFIO/n394 ), .A(pktrscendh) );
    snl_aoi033x0 \SAEXE/RFIO/U278  ( .ZN(\SAEXE/RFIO/n378 ), .A(pgadrovfh), 
        .B(\SAEXE/RFIO/fst[1] ), .C(\SAEXE/RFIO/fst[2] ), .D(
        \SAEXE/RFIO/phrefendh ), .E(\SAEXE/wrd_datah ), .F(
        \SAEXE/RFIO/phadrovfh ) );
    snl_aoi112x0 \SAEXE/RFIO/U236  ( .ZN(\SAEXE/RFIO/cnt4dech ), .A(
        \SAEXE/RFIO/n359 ), .B(\SAEXE/RFIO/n375 ), .C(\SAEXE/RFIO/n364 ), .D(
        pgadrovfh) );
    snl_nor02x1 \SAEXE/RFIO/U243  ( .ZN(ph_tbllt_h), .A(\SAEXE/RFIO/n386 ), 
        .B(\SAEXE/RFIO/n352 ) );
    snl_invx05 \SAEXE/RFIO/U258  ( .ZN(\SAEXE/RFIO/n353 ), .A(
        \SAEXE/RFIO/fst[0] ) );
    snl_nor02x1 \SAEXE/RFIO/U264  ( .ZN(\SAEXE/RFIO/n390 ), .A(
        \SAEXE/RFIO/n394 ), .B(\SAEXE/RFIO/n382 ) );
    snl_aoi022x1 \SAEXE/RFIO/U251  ( .ZN(\SAEXE/RFIO/n361 ), .A(
        \SAEXE/RFIO/n399 ), .B(\SAEXE/RFIO/n377 ), .C(\SAEXE/RFIO/n400 ), .D(
        \SAEXE/RFIO/n376 ) );
    snl_invx05 \SAEXE/RFIO/U276  ( .ZN(\SAEXE/RFIO/n388 ), .A(pktblcovfh) );
    snl_nor02x1 \SAEXE/RFIO/U281  ( .ZN(\SAEXE/RFIO/n406 ), .A(pktrscendh), 
        .B(\SAEXE/RFIO/cnt4out[3] ) );
    snl_nand13x1 \SAEXE/RFIO/U293  ( .ZN(\SAEXE/RFIO/n374 ), .A(pktblcendh), 
        .B(\SAEXE/RFIO/n390 ), .C(\SAEXE/RFIO/n389 ) );
    snl_invx05 \SAEXE/RFIO/U303  ( .ZN(\SAEXE/RFIO/n408 ), .A(\pk_psae_h[5] )
         );
    snl_invx1 \SAEXE/RFIO/U225  ( .ZN(\SAEXE/RFIO/n352 ), .A(\SAEXE/RFIO/n395 
        ) );
    snl_oai013x0 \SAEXE/RFIO/U237  ( .ZN(\SAEXE/adovflth2 ), .A(
        \SAEXE/RFIO/n376 ), .B(\SAEXE/RFIO/n377 ), .C(\SAEXE/RFIO/n353 ), .D(
        \SAEXE/RFIO/n378 ) );
    snl_nor02x1 \SAEXE/RFIO/U242  ( .ZN(ph_trscdech), .A(\SAEXE/RFIO/n385 ), 
        .B(\SAEXE/RFIO/n382 ) );
    snl_nor03x0 \SAEXE/RFIO/U265  ( .ZN(\SAEXE/RFIO/n389 ), .A(
        \SAEXE/RFIO/n360 ), .B(\SAEXE/RFIO/cnt4out[3] ), .C(\SAEXE/RFIO/n381 )
         );
    snl_nor02x1 \SAEXE/RFIO/U280  ( .ZN(\SAEXE/RFIO/n403 ), .A(pktblcendh), 
        .B(pktblcovfh) );
    snl_nand02x1 \SAEXE/RFIO/U288  ( .ZN(\SAEXE/RFIO/n356 ), .A(
        \SAEXE/RFIO/n389 ), .B(\SAEXE/RFIO/n407 ) );
    snl_ffqrnx1 \SAEXE/RFIO/fst_reg[3]  ( .Q(\SAEXE/trsc2_h ), .D(
        \SAEXE/RFIO/nfst[3] ), .RN(n10735), .CP(SCLK) );
    snl_nor02x1 \SAEXE/RFIO/U259  ( .ZN(\SAEXE/RFIO/*cell*3735/U62/CONTROL2 ), 
        .A(\SAEXE/RFIO/n353 ), .B(\SAEXE/RFIO/n357 ) );
    snl_oai223x0 \SAEXE/RFIO/U230  ( .ZN(\SAEXE/RFIO/nfst[2] ), .A(
        \SAEXE/RFIO/n357 ), .B(\SAEXE/RFIO/fst[0] ), .C(\SAEXE/RFIO/n358 ), 
        .D(\SAEXE/RFIO/n359 ), .E(\SAEXE/RFIO/n360 ), .F(\SAEXE/RFIO/n361 ), 
        .G(\SAEXE/RFIO/n362 ) );
    snl_nor02x1 \SAEXE/RFIO/U239  ( .ZN(ph_tblcdech), .A(pktblcendh), .B(
        \SAEXE/RFIO/n380 ) );
    snl_nor02x1 \SAEXE/RFIO/U250  ( .ZN(\SAEXE/RFIO/n358 ), .A(
        \SAEXE/RFIO/n398 ), .B(\SAEXE/RFIO/n366 ) );
    snl_invx05 \SAEXE/RFIO/U277  ( .ZN(\SAEXE/RFIO/n366 ), .A(ph_lberr) );
    snl_invx05 \SAEXE/RFIO/U289  ( .ZN(\SAEXE/RFIO/phrfin1h ), .A(
        \SAEXE/RFIO/n356 ) );
    snl_nand04x0 \SAEXE/RFIO/U292  ( .ZN(\SAEXE/RFIO/n402 ), .A(pktrscovfh), 
        .B(\SAEXE/RFIO/rfio1h ), .C(\SAEXE/RFIO/n406 ), .D(
        \SAEXE/RFIO/cnt4out[0] ) );
    snl_nand02x1 \SAEXE/RFIO/U302  ( .ZN(\SAEXE/RFIO/n375 ), .A(
        \SAEXE/RFIO/n407 ), .B(\SAEXE/RFIO/n386 ) );
    snl_oai012x1 \SAEXE/RFIO/U295  ( .ZN(\SAEXE/RFIO/n407 ), .A(pktrscendh), 
        .B(pktrscovfh), .C(\SAEXE/RFIO/rfio1h ) );
    snl_nand02x1 \SAEXE/RFIO/U257  ( .ZN(\SAEXE/RFIO/n357 ), .A(
        \SAEXE/RFIO/fst[2] ), .B(\SAEXE/RFIO/n362 ) );
    snl_nand03x0 \SAEXE/RFIO/U270  ( .ZN(\SAEXE/RFIO/n371 ), .A(
        \SAEXE/RFIO/n395 ), .B(\SAEXE/RFIO/rfio1h ), .C(\pk_psae_h[5] ) );
    snl_aoi012x1 \SAEXE/RFIO/U245  ( .ZN(\SAEXE/RFIO/n391 ), .A(pktblcendh), 
        .B(\SAEXE/RFIO/n353 ), .C(\SAEXE/RFIO/n362 ) );
    snl_nand04x0 \SAEXE/RFIO/U279  ( .ZN(\SAEXE/RFIO/n372 ), .A(\pk_psae_h[7] 
        ), .B(ph_saexe_sth), .C(\SAEXE/RFIO/n362 ), .D(\SAEXE/RFIO/n377 ) );
    snl_ffqrnx1 \SAEXE/RFIO/fst_reg[1]  ( .Q(\SAEXE/RFIO/fst[1] ), .D(
        \SAEXE/RFIO/nfst[1] ), .RN(n10735), .CP(SCLK) );
    snl_nor03x0 \SAEXE/RFIO/U262  ( .ZN(\SAEXE/RFIO/rfio1h ), .A(
        \SAEXE/RFIO/n404 ), .B(\pk_psae_h[6] ), .C(\pk_psae_h[4] ) );
    snl_invx05 \SAEXE/RFIO/U287  ( .ZN(\SAEXE/RFIO/n364 ), .A(
        \SAEXE/RFIO/*cell*3735/U62/CONTROL2 ) );
    snl_oai122x2 \SAEXE/RFIO/U227  ( .ZN(\SAEXE/RFIO/nfst[0] ), .A(ph_lberr), 
        .B(\SAEXE/RFIO/n352 ), .C(\SAEXE/RFIO/fst[2] ), .D(\SAEXE/RFIO/n353 ), 
        .E(\SAEXE/RFIO/n354 ) );
    snl_oai012x1 \SAEXE/RFIO/U229  ( .ZN(\SAEXE/RFIO/nfst[1] ), .A(
        \SAEXE/RFIO/fst[2] ), .B(\SAEXE/RFIO/n355 ), .C(\SAEXE/RFIO/n356 ) );
    snl_invx05 \SAEXE/RFIO/U255  ( .ZN(\SAEXE/RFIO/n362 ), .A(
        \SAEXE/RFIO/fst[1] ) );
    snl_invx05 \SAEXE/RFIO/U269  ( .ZN(\SAEXE/RFIO/n370 ), .A(
        \SAEXE/RFIO/cnt4out[1] ) );
    snl_nor03x0 \SAEXE/RFIO/U272  ( .ZN(\SAEXE/wrd_datah ), .A(
        \SAEXE/RFIO/fst[0] ), .B(\SAEXE/RFIO/fst[2] ), .C(\SAEXE/RFIO/n362 )
         );
    snl_ffqrnx1 \SAEXE/RFIO/fst_reg[0]  ( .Q(\SAEXE/RFIO/fst[0] ), .D(
        \SAEXE/RFIO/nfst[0] ), .RN(n10735), .CP(SCLK) );
    snl_invx05 \SAEXE/RFIO/U285  ( .ZN(\SAEXE/RFIO/n382 ), .A(
        \SAEXE/RFIO/rfio1h ) );
    snl_aoi012x1 \SAEXE/RFIO/U297  ( .ZN(\SAEXE/RFIO/n369 ), .A(
        \SAEXE/RFIO/n408 ), .B(\SAEXE/RFIO/rfio1h ), .C(\SAEXE/RFIO/rfin2h )
         );
    snl_oai023x0 \SAEXE/RFIO/U232  ( .ZN(ph_sa1lt_h), .A(\SAEXE/RFIO/n368 ), 
        .B(\SAEXE/RFIO/n369 ), .C(\SAEXE/RFIO/n352 ), .D(\SAEXE/RFIO/n370 ), 
        .E(\SAEXE/RFIO/n371 ) );
    snl_aoi013x0 \SAEXE/RFIO/U247  ( .ZN(\SAEXE/RFIO/n385 ), .A(
        \SAEXE/RFIO/n393 ), .B(\SAEXE/RFIO/n394 ), .C(\SAEXE/RFIO/n389 ), .D(
        \SAEXE/RFIO/ri1_trscdech ) );
    snl_nor02x1 \SAEXE/RFIO/U260  ( .ZN(\SAEXE/RFIO/n387 ), .A(
        \SAEXE/RFIO/n364 ), .B(pgadrovfh) );
    snl_nand12x1 \SAEXE/RFIO/U235  ( .ZN(\SAEXE/RFIO/reloadh ), .A(
        \SAEXE/RFIO/n373 ), .B(\SAEXE/RFIO/n374 ) );
    snl_nand12x1 \SAEXE/RFIO/U240  ( .ZN(\SAEXE/rf_srcadr1_h ), .A(
        \SAEXE/RFIO/srcadr1_h ), .B(\SAEXE/RFIO/n381 ) );
    snl_oai012x1 \SAEXE/RFIO/U299  ( .ZN(\SAEXE/RFIO/n400 ), .A(pktblcendh), 
        .B(\SAEXE/RFIO/n377 ), .C(\SAEXE/RFIO/n353 ) );
    snl_aoi122x0 \SAEXE/RFIO/U249  ( .ZN(\SAEXE/RFIO/n363 ), .A(pktblcendh), 
        .B(\SAEXE/RFIO/n396 ), .C(pktblcovfh), .D(\SAEXE/RFIO/cnt4out[3] ), 
        .E(\SAEXE/RFIO/n397 ) );
    snl_aoi012x1 \SAEXE/RFIO/U252  ( .ZN(\SAEXE/RFIO/n355 ), .A(
        \SAEXE/RFIO/fst[1] ), .B(\SAEXE/RFIO/n401 ), .C(\SAEXE/RFIO/fst[0] )
         );
    snl_invx05 \SAEXE/RFIO/U267  ( .ZN(\SAEXE/RFIO/n398 ), .A(ph_lbend) );
    snl_nand02x1 \SAEXE/RFIO/U282  ( .ZN(\SAEXE/RFIO/n397 ), .A(
        \SAEXE/RFIO/n402 ), .B(\SAEXE/RFIO/n376 ) );
    snl_oai112x0 \SAEXE/RFIO/U290  ( .ZN(\SAEXE/RFIO/n384 ), .A(
        \SAEXE/RFIO/n391 ), .B(\SAEXE/RFIO/n392 ), .C(\SAEXE/RFIO/n376 ), .D(
        \SAEXE/RFIO/fst[2] ) );
    snl_oai013x0 \SAEXE/RFIO/U300  ( .ZN(\SAEXE/RFIO/n399 ), .A(
        \SAEXE/RFIO/n405 ), .B(ph_lberr), .C(\SAEXE/RFIO/phadrovfh ), .D(
        \SAEXE/RFIO/n353 ) );
    snl_ffqrnx1 \SAEXE/RFIO/fst_reg[2]  ( .Q(\SAEXE/RFIO/fst[2] ), .D(
        \SAEXE/RFIO/nfst[2] ), .RN(n10735), .CP(SCLK) );
    snl_invx05 \SAEXE/RFIO/U275  ( .ZN(\SAEXE/RFIO/n393 ), .A(pktrscovfh) );
    snl_nand12x1 \SAEXE/RFIO/U226  ( .ZN(\SAEXE/n434 ), .A(
        \SAEXE/RFIO/RIN1TRS ), .B(\SAEXE/RFIO/n383 ) );
    snl_ao01b2x0 \SAEXE/RFIO/U234  ( .Z(\SAEXE/RFIO/cntloadh ), .A(
        \SAEXE/RFIO/fst[0] ), .B(\SAEXE/RFIO/n372 ), .C(\SAEXE/trsc2_h ) );
    snl_nand12x1 \SAEXE/RFIO/U241  ( .ZN(\SAEXE/sa_start3 ), .A(
        \SAEXE/RFIO/phrfin1sah ), .B(\SAEXE/RFIO/n384 ) );
    snl_aoi0b12x0 \SAEXE/RFIO/U283  ( .ZN(\SAEXE/RFIO/n367 ), .A(pktblcendh), 
        .B(\SAEXE/RFIO/n373 ), .C(\SAEXE/RFIO/n378 ) );
    snl_ffqx1 \SAEXE/RFIO/RIN1TRS_reg  ( .Q(\SAEXE/RFIO/RIN1TRS ), .D(
        \SAEXE/RFIO/rfin1tpenh ), .CP(SCLK) );
    snl_nor03x0 \SAEXE/RFIO/U266  ( .ZN(\SAEXE/RFIO/n373 ), .A(
        \SAEXE/RFIO/n362 ), .B(\SAEXE/RFIO/fst[0] ), .C(\SAEXE/RFIO/n377 ) );
    snl_ao012x1 \SAEXE/RFIO/U298  ( .Z(\SAEXE/RFIO/n396 ), .A(
        \SAEXE/RFIO/cnt4out[0] ), .B(\SAEXE/RFIO/n390 ), .C(
        \SAEXE/RFIO/cnt4out[3] ) );
    snl_nor03x1 \SAEXE/RFIO/U228  ( .ZN(ph_trslt_h), .A(\SAEXE/RFIO/n352 ), 
        .B(\SAEXE/RFIO/n381 ), .C(\SAEXE/RFIO/n382 ) );
    snl_oai023x0 \SAEXE/RFIO/U233  ( .ZN(ph_sa2lt_h), .A(\SAEXE/RFIO/n370 ), 
        .B(\SAEXE/RFIO/n369 ), .C(\SAEXE/RFIO/n352 ), .D(\SAEXE/RFIO/n371 ), 
        .E(\SAEXE/RFIO/n368 ) );
    snl_aoi012x1 \SAEXE/RFIO/U248  ( .ZN(\SAEXE/RFIO/n365 ), .A(
        \SAEXE/RFIO/phrefendh ), .B(\SAEXE/wrd_datah ), .C(\SAEXE/RFIO/n395 )
         );
    snl_oa013x1 \SAEXE/RFIO/U253  ( .Z(\SAEXE/RFIO/n379 ), .A(
        \SAEXE/RFIO/n386 ), .B(pktblcendh), .C(\SAEXE/RFIO/n388 ), .D(
        \SAEXE/RFIO/n402 ) );
    snl_aoi022x1 \SAEXE/RFIO/U254  ( .ZN(\SAEXE/RFIO/n359 ), .A(
        \SAEXE/RFIO/n403 ), .B(\SAEXE/RFIO/cnt4out[3] ), .C(\SAEXE/RFIO/n381 ), 
        .D(\SAEXE/RFIO/n386 ) );
    snl_invx05 \SAEXE/RFIO/U273  ( .ZN(\SAEXE/RFIO/n405 ), .A(
        \SAEXE/RFIO/phrefendh ) );
    snl_invx05 \SAEXE/RFIO/U274  ( .ZN(\SAEXE/RFIO/n376 ), .A(pgadrovfh) );
    snl_invx05 \SAEXE/RFIO/U291  ( .ZN(ph_tpralt_h), .A(\SAEXE/RFIO/n384 ) );
    snl_oai012x1 \SAEXE/RFIO/U296  ( .ZN(\SAEXE/RFIO/n383 ), .A(
        \SAEXE/RFIO/fst[0] ), .B(\SAEXE/RFIO/fst[2] ), .C(\SAEXE/RFIO/n381 )
         );
    snl_oai012x1 \SAEXE/RFIO/U301  ( .ZN(\SAEXE/RFIO/n401 ), .A(ph_lberr), .B(
        \SAEXE/RFIO/phadrovfh ), .C(\SAEXE/RFIO/phrefendh ) );
    snl_nor03x0 \SAEXE/RFIO/U268  ( .ZN(\SAEXE/RFIO/n395 ), .A(
        \SAEXE/RFIO/n357 ), .B(\SAEXE/RFIO/fst[0] ), .C(\SAEXE/RFIO/n398 ) );
    snl_nor02x1 \SAEXE/RFIO/U246  ( .ZN(\SAEXE/RFIO/n392 ), .A(
        \SAEXE/RFIO/n359 ), .B(\SAEXE/RFIO/n353 ) );
    snl_invx05 \SAEXE/RFIO/U261  ( .ZN(\SAEXE/RFIO/n381 ), .A(
        \SAEXE/RFIO/cnt4out[0] ) );
    snl_oa012x1 \SAEXE/RFIO/U284  ( .Z(\SAEXE/RFIO/n354 ), .A(
        \SAEXE/RFIO/n372 ), .B(\SAEXE/trsc2_h ), .C(\SAEXE/RFIO/n374 ) );
    snl_sffqrnx1 \SAEXE/RFIO/ph_tcer_h_reg  ( .Q(ph_tcer_h), .D(1'b0), .RN(
        n10735), .SD(\SAEXE/RFIO/*cell*3735/U62/CONTROL2 ), .SE(
        \SAEXE/RFIO/*cell*3735/U61/Z_0 ), .CP(SCLK) );
    snl_bufx1 \SADR/SELOPR/U8  ( .Z(\SADR/SELOPR/n10656 ), .A(ph_tprsel_h) );
    snl_nand02x1 \SADR/SELOPR/U13  ( .ZN(\SADR/operand[23] ), .A(
        \SADR/SELOPR/n10665 ), .B(\SADR/SELOPR/n10666 ) );
    snl_nand02x1 \SADR/SELOPR/U14  ( .ZN(\SADR/operand[22] ), .A(
        \SADR/SELOPR/n10667 ), .B(\SADR/SELOPR/n10668 ) );
    snl_nand02x1 \SADR/SELOPR/U21  ( .ZN(\SADR/operand[15] ), .A(
        \SADR/SELOPR/n10681 ), .B(\SADR/SELOPR/n10682 ) );
    snl_aoi222x0 \SADR/SELOPR/U54  ( .ZN(\SADR/SELOPR/n10695 ), .A(
        \pk_trba_h[8] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[8] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[8] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U73  ( .ZN(\SADR/SELOPR/n10730 ), .A(
        \pk_dpr_h[28] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[28] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[28] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U113  ( .ZN(\SADR/SELOPR/n10712 ), .A(
        \pk_dpr_h[0] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[0] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[0] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U96  ( .ZN(\SADR/SELOPR/n10675 ), .A(
        \pk_trba_h[18] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[18] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[18] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U68  ( .ZN(\SADR/SELOPR/n10723 ), .A(
        \pk_trba_h[30] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[30] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[30] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U108  ( .ZN(\SADR/SELOPR/n10687 ), .A(
        \pk_trba_h[12] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[12] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[12] ), .F(\SADR/SELOPR/n10718 ) );
    snl_nand02x1 \SADR/SELOPR/U28  ( .ZN(\SADR/operand[8] ), .A(
        \SADR/SELOPR/n10695 ), .B(\SADR/SELOPR/n10696 ) );
    snl_nand02x1 \SADR/SELOPR/U33  ( .ZN(\SADR/operand[3] ), .A(
        \SADR/SELOPR/n10705 ), .B(\SADR/SELOPR/n10706 ) );
    snl_nand02x1 \SADR/SELOPR/U34  ( .ZN(\SADR/operand[2] ), .A(
        \SADR/SELOPR/n10707 ), .B(\SADR/SELOPR/n10708 ) );
    snl_and02x1 \SADR/SELOPR/U41  ( .Z(\SADR/SELOPR/n10718 ), .A(ph_oprtrs_h), 
        .B(\SADR/SELOPR/n10714 ) );
    snl_mux21x1 \SADR/SELOPR/U46  ( .Z(\pgsdprhh[30] ), .A(
        \SADR/SELOPR/n10722 ), .B(\SADR/m_fadrh[30] ), .S(pgfbadrsel) );
    snl_aoi222x0 \SADR/SELOPR/U61  ( .ZN(\SADR/SELOPR/n10704 ), .A(
        \pk_dpr_h[4] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[4] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[4] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U84  ( .ZN(\SADR/SELOPR/n10665 ), .A(
        \pk_trba_h[23] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[23] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[23] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U101  ( .ZN(\SADR/SELOPR/n10682 ), .A(
        \pk_dpr_h[15] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[15] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[15] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U66  ( .ZN(\SADR/SELOPR/n10720 ), .A(
        \pk_trba_h[31] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[31] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[31] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U106  ( .ZN(\SADR/SELOPR/n10685 ), .A(
        \pk_trba_h[13] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[13] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[13] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U83  ( .ZN(\SADR/SELOPR/n10666 ), .A(
        \pk_dpr_h[23] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[23] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[23] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U98  ( .ZN(\SADR/SELOPR/n10677 ), .A(
        \pk_trba_h[17] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[17] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[17] ), .F(\SADR/SELOPR/n10718 ) );
    snl_nand02x1 \SADR/SELOPR/U26  ( .ZN(\SADR/operand[10] ), .A(
        \SADR/SELOPR/n10691 ), .B(\SADR/SELOPR/n10692 ) );
    snl_mux21x1 \SADR/SELOPR/U48  ( .Z(\pgsdprhh[29] ), .A(
        \SADR/SELOPR/n10725 ), .B(\SADR/m_fadrh[29] ), .S(pgfbadrsel) );
    snl_nand02x1 \SADR/SELOPR/U9  ( .ZN(\SADR/operand[27] ), .A(
        \SADR/SELOPR/n10657 ), .B(\SADR/SELOPR/n10658 ) );
    snl_nand02x1 \SADR/SELOPR/U12  ( .ZN(\SADR/operand[24] ), .A(
        \SADR/SELOPR/n10663 ), .B(\SADR/SELOPR/n10664 ) );
    snl_nand02x1 \SADR/SELOPR/U35  ( .ZN(\SADR/operand[1] ), .A(
        \SADR/SELOPR/n10709 ), .B(\SADR/SELOPR/n10710 ) );
    snl_aoi222x0 \SADR/SELOPR/U53  ( .ZN(\SADR/SELOPR/n10696 ), .A(
        \pk_dpr_h[8] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[8] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[8] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U91  ( .ZN(\SADR/SELOPR/n10710 ), .A(
        \pk_dpr_h[1] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[1] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[1] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U74  ( .ZN(\SADR/SELOPR/n10729 ), .A(
        \pk_trba_h[28] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[28] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[28] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U114  ( .ZN(\SADR/SELOPR/n10711 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(\pk_spr_h[0] ), .D(\SADR/SELOPR/n10717 ), 
        .E(\stream3[0] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U99  ( .ZN(\SADR/SELOPR/n10680 ), .A(
        \pk_dpr_h[16] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[16] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[16] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_nand02x1 \SADR/SELOPR/U27  ( .ZN(\SADR/operand[9] ), .A(
        \SADR/SELOPR/n10693 ), .B(\SADR/SELOPR/n10694 ) );
    snl_and12x1 \SADR/SELOPR/U40  ( .Z(\SADR/SELOPR/n10717 ), .A(
        \SADR/SELOPR/n10656 ), .B(ph_sprtrs_h) );
    snl_aoi222x0 \SADR/SELOPR/U82  ( .ZN(\SADR/SELOPR/n10663 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(1'b0), .D(\SADR/SELOPR/n10717 ), .E(
        \stream3[24] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U52  ( .ZN(\SADR/SELOPR/n10693 ), .A(
        \SADR/SELOPR/n10656 ), .B(\pk_trba_h[9] ), .C(\pk_spr_h[9] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[9] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U67  ( .ZN(\SADR/SELOPR/n10724 ), .A(
        \pk_dpr_h[30] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[30] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[30] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U107  ( .ZN(\SADR/SELOPR/n10688 ), .A(
        \pk_dpr_h[12] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[12] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[12] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U75  ( .ZN(\SADR/SELOPR/n10658 ), .A(1'b0), .B(
        \SADR/SELOPR/n10716 ), .C(1'b0), .D(\SADR/SELOPR/n10713 ), .E(1'b0), 
        .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U90  ( .ZN(\SADR/SELOPR/n10671 ), .A(
        \pk_trba_h[20] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[20] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[20] ), .F(\SADR/SELOPR/n10718 ) );
    snl_nand02x1 \SADR/SELOPR/U10  ( .ZN(\SADR/operand[26] ), .A(
        \SADR/SELOPR/n10659 ), .B(\SADR/SELOPR/n10660 ) );
    snl_nand02x1 \SADR/SELOPR/U15  ( .ZN(\SADR/operand[21] ), .A(
        \SADR/SELOPR/n10669 ), .B(\SADR/SELOPR/n10670 ) );
    snl_nand02x1 \SADR/SELOPR/U20  ( .ZN(\SADR/operand[16] ), .A(
        \SADR/SELOPR/n10679 ), .B(\SADR/SELOPR/n10680 ) );
    snl_nand02x1 \SADR/SELOPR/U49  ( .ZN(\SADR/SELOPR/n10728 ), .A(
        \SADR/SELOPR/n10729 ), .B(\SADR/SELOPR/n10730 ) );
    snl_aoi222x0 \SADR/SELOPR/U69  ( .ZN(\SADR/SELOPR/n10708 ), .A(
        \pk_dpr_h[2] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[2] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[2] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U109  ( .ZN(\SADR/SELOPR/n10690 ), .A(
        \pk_dpr_h[11] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[11] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[11] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_nand02x1 \SADR/SELOPR/U29  ( .ZN(\SADR/operand[7] ), .A(
        \SADR/SELOPR/n10697 ), .B(\SADR/SELOPR/n10698 ) );
    snl_nand02x1 \SADR/SELOPR/U47  ( .ZN(\SADR/SELOPR/n10725 ), .A(
        \SADR/SELOPR/n10726 ), .B(\SADR/SELOPR/n10727 ) );
    snl_aoi222x0 \SADR/SELOPR/U55  ( .ZN(\SADR/SELOPR/n10698 ), .A(
        \pk_dpr_h[7] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[7] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[7] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U72  ( .ZN(\SADR/SELOPR/n10726 ), .A(
        \pk_trba_h[29] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[29] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[29] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U97  ( .ZN(\SADR/SELOPR/n10678 ), .A(
        \pk_dpr_h[17] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[17] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[17] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U112  ( .ZN(\SADR/SELOPR/n10691 ), .A(
        \pk_trba_h[10] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[10] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[10] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U60  ( .ZN(\SADR/SELOPR/n10701 ), .A(
        \pk_trba_h[5] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[5] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[5] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U100  ( .ZN(\SADR/SELOPR/n10679 ), .A(
        \pk_trba_h[16] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[16] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[16] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U85  ( .ZN(\SADR/SELOPR/n10668 ), .A(
        \pk_dpr_h[22] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[22] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[22] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_nand02x1 \SADR/SELOPR/U17  ( .ZN(\SADR/operand[19] ), .A(
        \SADR/SELOPR/n10673 ), .B(\SADR/SELOPR/n10674 ) );
    snl_nand02x1 \SADR/SELOPR/U22  ( .ZN(\SADR/operand[14] ), .A(
        \SADR/SELOPR/n10683 ), .B(\SADR/SELOPR/n10684 ) );
    snl_nand02x1 \SADR/SELOPR/U32  ( .ZN(\SADR/operand[4] ), .A(
        \SADR/SELOPR/n10703 ), .B(\SADR/SELOPR/n10704 ) );
    snl_and02x1 \SADR/SELOPR/U39  ( .Z(\SADR/SELOPR/n10716 ), .A(ph_dprtrs_h), 
        .B(\SADR/SELOPR/n10714 ) );
    snl_aoi222x0 \SADR/SELOPR/U57  ( .ZN(\SADR/SELOPR/n10700 ), .A(
        \pk_dpr_h[6] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[6] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[6] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U70  ( .ZN(\SADR/SELOPR/n10707 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(\pk_spr_h[2] ), .D(\SADR/SELOPR/n10717 ), 
        .E(\stream3[2] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U110  ( .ZN(\SADR/SELOPR/n10689 ), .A(
        \pk_trba_h[11] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[11] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[11] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U95  ( .ZN(\SADR/SELOPR/n10676 ), .A(
        \pk_dpr_h[18] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[18] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[18] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_nand02x1 \SADR/SELOPR/U30  ( .ZN(\SADR/operand[6] ), .A(
        \SADR/SELOPR/n10699 ), .B(\SADR/SELOPR/n10700 ) );
    snl_aoi222x0 \SADR/SELOPR/U79  ( .ZN(\SADR/SELOPR/n10662 ), .A(1'b0), .B(
        \SADR/SELOPR/n10716 ), .C(1'b0), .D(\SADR/SELOPR/n10713 ), .E(1'b0), 
        .F(\SADR/SELOPR/n10715 ) );
    snl_invx05 \SADR/SELOPR/U42  ( .ZN(\SADR/SELOPR/n10714 ), .A(
        \SADR/SELOPR/n10656 ) );
    snl_nand02x1 \SADR/SELOPR/U45  ( .ZN(\SADR/SELOPR/n10722 ), .A(
        \SADR/SELOPR/n10723 ), .B(\SADR/SELOPR/n10724 ) );
    snl_aoi222x0 \SADR/SELOPR/U87  ( .ZN(\SADR/SELOPR/n10670 ), .A(
        \pk_dpr_h[21] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[21] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[21] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U62  ( .ZN(\SADR/SELOPR/n10703 ), .A(
        \pk_trba_h[4] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[4] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[4] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U65  ( .ZN(\SADR/SELOPR/n10721 ), .A(
        \pk_dpr_h[31] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[31] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[31] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U102  ( .ZN(\SADR/SELOPR/n10681 ), .A(
        \pk_trba_h[15] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[15] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[15] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U105  ( .ZN(\SADR/SELOPR/n10686 ), .A(
        \pk_dpr_h[13] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[13] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[13] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U80  ( .ZN(\SADR/SELOPR/n10661 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(1'b0), .D(\SADR/SELOPR/n10717 ), .E(
        \stream3[25] ), .F(\SADR/SELOPR/n10718 ) );
    snl_nand02x1 \SADR/SELOPR/U11  ( .ZN(\SADR/operand[25] ), .A(
        \SADR/SELOPR/n10661 ), .B(\SADR/SELOPR/n10662 ) );
    snl_nand02x1 \SADR/SELOPR/U19  ( .ZN(\SADR/operand[17] ), .A(
        \SADR/SELOPR/n10677 ), .B(\SADR/SELOPR/n10678 ) );
    snl_nand02x1 \SADR/SELOPR/U25  ( .ZN(\SADR/operand[11] ), .A(
        \SADR/SELOPR/n10689 ), .B(\SADR/SELOPR/n10690 ) );
    snl_and02x1 \SADR/SELOPR/U37  ( .Z(\SADR/SELOPR/n10713 ), .A(ph_srcadr2_h), 
        .B(\SADR/SELOPR/n10714 ) );
    snl_aoi222x0 \SADR/SELOPR/U59  ( .ZN(\SADR/SELOPR/n10702 ), .A(
        \pk_dpr_h[5] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[5] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[5] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U89  ( .ZN(\SADR/SELOPR/n10672 ), .A(
        \pk_dpr_h[20] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[20] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[20] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_mux21x1 \SADR/SELOPR/U50  ( .Z(\pgsdprhh[28] ), .A(
        \SADR/SELOPR/n10728 ), .B(\SADR/m_fadrh[28] ), .S(pgfbadrsel) );
    snl_aoi222x0 \SADR/SELOPR/U77  ( .ZN(\SADR/SELOPR/n10660 ), .A(1'b0), .B(
        \SADR/SELOPR/n10716 ), .C(1'b0), .D(\SADR/SELOPR/n10713 ), .E(1'b0), 
        .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U92  ( .ZN(\SADR/SELOPR/n10709 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(\pk_spr_h[1] ), .D(\SADR/SELOPR/n10717 ), 
        .E(\stream3[1] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U58  ( .ZN(\SADR/SELOPR/n10699 ), .A(
        \pk_trba_h[6] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[6] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[6] ), .F(\SADR/SELOPR/n10718 ) );
    snl_nand02x1 \SADR/SELOPR/U16  ( .ZN(\SADR/operand[20] ), .A(
        \SADR/SELOPR/n10671 ), .B(\SADR/SELOPR/n10672 ) );
    snl_nand02x1 \SADR/SELOPR/U18  ( .ZN(\SADR/operand[18] ), .A(
        \SADR/SELOPR/n10675 ), .B(\SADR/SELOPR/n10676 ) );
    snl_nand02x1 \SADR/SELOPR/U36  ( .ZN(\SADR/operand[0] ), .A(
        \SADR/SELOPR/n10711 ), .B(\SADR/SELOPR/n10712 ) );
    snl_nand02x1 \SADR/SELOPR/U43  ( .ZN(\SADR/SELOPR/n10719 ), .A(
        \SADR/SELOPR/n10720 ), .B(\SADR/SELOPR/n10721 ) );
    snl_aoi222x0 \SADR/SELOPR/U64  ( .ZN(\SADR/SELOPR/n10705 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(\pk_spr_h[3] ), .D(\SADR/SELOPR/n10717 ), 
        .E(\stream3[3] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U81  ( .ZN(\SADR/SELOPR/n10664 ), .A(1'b0), .B(
        \SADR/SELOPR/n10716 ), .C(1'b0), .D(\SADR/SELOPR/n10713 ), .E(1'b0), 
        .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U104  ( .ZN(\SADR/SELOPR/n10683 ), .A(
        \pk_trba_h[14] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[14] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[14] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U51  ( .ZN(\SADR/SELOPR/n10694 ), .A(
        \pk_dpr_h[9] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[9] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[9] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U76  ( .ZN(\SADR/SELOPR/n10657 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(1'b0), .D(\SADR/SELOPR/n10717 ), .E(
        \stream3[27] ), .F(\SADR/SELOPR/n10718 ) );
    snl_nand02x1 \SADR/SELOPR/U23  ( .ZN(\SADR/operand[13] ), .A(
        \SADR/SELOPR/n10685 ), .B(\SADR/SELOPR/n10686 ) );
    snl_nand02x1 \SADR/SELOPR/U24  ( .ZN(\SADR/operand[12] ), .A(
        \SADR/SELOPR/n10687 ), .B(\SADR/SELOPR/n10688 ) );
    snl_aoi222x0 \SADR/SELOPR/U88  ( .ZN(\SADR/SELOPR/n10669 ), .A(
        \pk_trba_h[21] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[21] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[21] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U93  ( .ZN(\SADR/SELOPR/n10674 ), .A(
        \pk_dpr_h[19] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[19] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[19] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_nand02x1 \SADR/SELOPR/U31  ( .ZN(\SADR/operand[5] ), .A(
        \SADR/SELOPR/n10701 ), .B(\SADR/SELOPR/n10702 ) );
    snl_and02x1 \SADR/SELOPR/U38  ( .Z(\SADR/SELOPR/n10715 ), .A(ph_srcadr1_h), 
        .B(\SADR/SELOPR/n10714 ) );
    snl_mux21x1 \SADR/SELOPR/U44  ( .Z(\pgsdprhh[31] ), .A(
        \SADR/SELOPR/n10719 ), .B(\SADR/m_fadrh[31] ), .S(pgfbadrsel) );
    snl_aoi222x0 \SADR/SELOPR/U56  ( .ZN(\SADR/SELOPR/n10697 ), .A(
        \pk_trba_h[7] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[7] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[7] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U94  ( .ZN(\SADR/SELOPR/n10673 ), .A(
        \pk_trba_h[19] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[19] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[19] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U71  ( .ZN(\SADR/SELOPR/n10727 ), .A(
        \pk_dpr_h[29] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[29] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[29] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U111  ( .ZN(\SADR/SELOPR/n10692 ), .A(
        \pk_dpr_h[10] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[10] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[10] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U63  ( .ZN(\SADR/SELOPR/n10706 ), .A(
        \pk_dpr_h[3] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[3] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[3] ), .F(\SADR/SELOPR/n10715 ) );
    snl_aoi222x0 \SADR/SELOPR/U86  ( .ZN(\SADR/SELOPR/n10667 ), .A(
        \pk_trba_h[22] ), .B(\SADR/SELOPR/n10656 ), .C(\pk_spr_h[22] ), .D(
        \SADR/SELOPR/n10717 ), .E(\stream3[22] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/SELOPR/U103  ( .ZN(\SADR/SELOPR/n10684 ), .A(
        \pk_dpr_h[14] ), .B(\SADR/SELOPR/n10716 ), .C(\pk_sra2_h[14] ), .D(
        \SADR/SELOPR/n10713 ), .E(\pk_sra1_h[14] ), .F(\SADR/SELOPR/n10715 )
         );
    snl_aoi222x0 \SADR/SELOPR/U78  ( .ZN(\SADR/SELOPR/n10659 ), .A(1'b0), .B(
        \SADR/SELOPR/n10656 ), .C(1'b0), .D(\SADR/SELOPR/n10717 ), .E(
        \stream3[26] ), .F(\SADR/SELOPR/n10718 ) );
    snl_aoi222x0 \SADR/MAINSADR/U14  ( .ZN(\SADR/MAINSADR/n8668 ), .A(
        \SADR/MAINSADR/oddadd_m1[23] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[22] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[22] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U21  ( .ZN(\SADR/MAINSADR/n8784 ), .A(
        \SADR/MAINSADR/oddadd_m1[16] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[15] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[15] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_nor02x1 \SADR/MAINSADR/U54  ( .ZN(\SADR/MAINSADR/offset[20] ), .A(
        \SADR/MAINSADR/n8643 ), .B(\SADR/MAINSADR/n8644 ) );
    snl_muxi21x1 \SADR/MAINSADR/U73  ( .ZN(\SADR/MAINSADR/n8681 ), .A(
        \SADR/MAINSADR/addindoff[10] ), .B(\SADR/m_fadrl[14] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_nor02x1 \SADR/MAINSADR/U113  ( .ZN(\SADR/MAINSADR/n8713 ), .A(
        \SADR/operand[26] ), .B(\SADR/operand[27] ) );
    snl_muxi21x1 \SADR/MAINSADR/U223  ( .ZN(\SADR/MAINSADR/index[18] ), .A(
        \SADR/MAINSADR/n8872 ), .B(\SADR/MAINSADR/n8877 ), .S(ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U432  ( .ZN(\SADR/MAINSADR/oddadd[13] ), .A(
        \SADR/MAINSADR/n8693 ) );
    snl_muxi21x1 \SADR/MAINSADR/U134  ( .ZN(\pgregadrh[9] ), .A(
        \SADR/MAINSADR/n8748 ), .B(\SADR/MAINSADR/n8745 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_nand03x0 \SADR/MAINSADR/U96  ( .ZN(\SADR/MAINSADR/n8663 ), .A(
        \SADR/MAINSADR/n8696 ), .B(ph_lwdsrc_h), .C(ph_adrdec_h) );
    snl_muxi21x1 \SADR/MAINSADR/U198  ( .ZN(\SADR/MAINSADR/index[9] ), .A(
        \SADR/MAINSADR/n8814 ), .B(\SADR/MAINSADR/n8819 ), .S(ph_lwdsrc_h) );
    snl_muxi21x1 \SADR/MAINSADR/U204  ( .ZN(\SADR/MAINSADR/index[6] ), .A(
        \SADR/MAINSADR/n8829 ), .B(\SADR/MAINSADR/n8834 ), .S(ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U394  ( .ZN(\SADR/MAINSADR/n8859 ), .A(
        \SADR/MAINSADR/n8725 ) );
    snl_muxi21x1 \SADR/MAINSADR/U415  ( .ZN(\pgsdprlh[7] ), .A(
        \SADR/MAINSADR/n8685 ), .B(\SADR/MAINSADR/n8678 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U338  ( .ZN(\SADR/MAINSADR/n8909 ), .A(
        \SADR/pgaddwz[11] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[11] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[11] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[11] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_nand02x1 \SADR/MAINSADR/U356  ( .ZN(\SADR/MAINSADR/n8648 ), .A(
        \SADR/MAINSADR/n8634 ), .B(\SADR/MAINSADR/oddadd[0] ) );
    snl_invx05 \SADR/MAINSADR/U371  ( .ZN(\SADR/MAINSADR/oddadd[20] ), .A(
        \SADR/MAINSADR/n8640 ) );
    snl_muxi21x1 \SADR/MAINSADR/U166  ( .ZN(\pgregadrh[16] ), .A(
        \SADR/MAINSADR/n8794 ), .B(\SADR/MAINSADR/n8782 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_nor03x0 \SADR/MAINSADR/U256  ( .ZN(\SADR/MAINSADR/n8919 ), .A(
        \SADR/MAINSADR/ovf_addindoff ), .B(\SADR/MAINSADR/oddadd[23] ), .C(
        \SADR/seglmterr ) );
    snl_aoi222x0 \SADR/MAINSADR/U271  ( .ZN(\SADR/MAINSADR/n8820 ), .A(
        \pk_indw_h[8] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[8] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[8] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U68  ( .ZN(\SADR/MAINSADR/n8675 ), .A(
        \SADR/MAINSADR/addindoff[8] ), .B(\SADR/m_fadrl[12] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U108  ( .Z(\SADR/MAINSADR/n8708 ), .A(
        \SADR/MAINSADR/n8707 ), .B(\SADR/MAINSADR/n8702 ) );
    snl_oa112x1 \SADR/MAINSADR/U141  ( .Z(\SADR/MAINSADR/n8763 ), .A(
        \SADR/MAINSADR/n8680 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8764 ), .D(\SADR/MAINSADR/n8765 ) );
    snl_muxi21x1 \SADR/MAINSADR/U183  ( .ZN(\SADR/MAINSADR/offset[2] ), .A(
        \SADR/MAINSADR/n8808 ), .B(\SADR/MAINSADR/n8651 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U294  ( .ZN(\SADR/MAINSADR/n8851 ), .A(
        \SADR/pgaddwz[2] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[2] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[2] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[2] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U304  ( .ZN(\SADR/MAINSADR/n8871 ), .A(
        \SADR/pgaddwxyz[0] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[0] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[0] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[0] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_aoi222x0 \SADR/MAINSADR/U323  ( .ZN(\SADR/MAINSADR/n8888 ), .A(
        \pk_indw_h[15] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[15] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[15] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U238  ( .ZN(\SADR/MAINSADR/index[10] ), .A(
        \SADR/MAINSADR/n8912 ), .B(\SADR/MAINSADR/n8814 ), .S(ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U429  ( .ZN(\SADR/MAINSADR/oddadd[15] ), .A(
        \SADR/MAINSADR/n8691 ) );
    snl_muxi21x1 \SADR/MAINSADR/U174  ( .ZN(\pgregadrh[10] ), .A(
        \SADR/MAINSADR/n8763 ), .B(\SADR/MAINSADR/n8800 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_muxi21x1 \SADR/MAINSADR/U191  ( .ZN(\SADR/MAINSADR/offset[13] ), .A(
        \SADR/MAINSADR/n8811 ), .B(\SADR/MAINSADR/n8803 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U286  ( .ZN(\SADR/MAINSADR/n8841 ), .A(
        \SADR/pgaddwz[4] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[4] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[4] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[4] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U316  ( .ZN(\SADR/MAINSADR/n8886 ), .A(
        \SADR/pgaddwxyz[16] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[16] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[16] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[16] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi222x0 \SADR/MAINSADR/U331  ( .ZN(\SADR/MAINSADR/n8898 ), .A(
        \pk_indw_h[13] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[13] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[13] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_nand02x1 \SADR/MAINSADR/U378  ( .ZN(\SADR/MAINSADR/n8758 ), .A(
        \SADR/MAINSADR/oddadd_p1[7] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U244  ( .ZN(\SADR/MAINSADR/n8734 ), .A(
        \SADR/pgaddwxyz[22] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[22] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[22] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[22] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi222x0 \SADR/MAINSADR/U28  ( .ZN(\SADR/MAINSADR/n8747 ), .A(
        \SADR/MAINSADR/n8698 ), .B(\SADR/MAINSADR/oddadd_m1[9] ), .C(
        \SADR/MAINSADR/n8917 ), .D(\SADR/MAINSADR/oddadd_m2[8] ), .E(
        \SADR/MAINSADR/n8918 ), .F(\SADR/MAINSADR/oddadd_p2[8] ) );
    snl_aoi222x0 \SADR/MAINSADR/U33  ( .ZN(\SADR/MAINSADR/n8750 ), .A(
        \SADR/MAINSADR/oddadd_m1[5] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[4] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[4] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_and05x1 \SADR/MAINSADR/U263  ( .Z(\SADR/MAINSADR/n8659 ), .A(
        \SADR/MAINSADR/cmpflg ), .B(\SADR/MAINSADR/n8928 ), .C(
        \SADR/MAINSADR/n8927 ), .D(\SADR/MAINSADR/n8926 ), .E(
        \SADR/MAINSADR/n8925 ) );
    snl_muxi21x1 \SADR/MAINSADR/U148  ( .ZN(\pgregadrh[3] ), .A(
        \SADR/MAINSADR/n8653 ), .B(\SADR/MAINSADR/n8760 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_muxi21x1 \SADR/MAINSADR/U153  ( .ZN(\pgregadrh[22] ), .A(
        \SADR/MAINSADR/n8776 ), .B(\SADR/MAINSADR/n8669 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x2 \SADR/MAINSADR/U41  ( .ZN(\pgsdprlh[15] ), .A(
        \SADR/MAINSADR/n8679 ), .B(\SADR/MAINSADR/n8691 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_invx1 \SADR/MAINSADR/U46  ( .ZN(\SADR/MAINSADR/n8917 ), .A(
        \SADR/MAINSADR/n8663 ) );
    snl_oai012x1 \SADR/MAINSADR/U61  ( .ZN(\pgsdprlh[3] ), .A(
        \SADR/MAINSADR/n8635 ), .B(\SADR/MAINSADR/n8653 ), .C(
        \SADR/MAINSADR/n8654 ) );
    snl_muxi21x1 \SADR/MAINSADR/U84  ( .ZN(\SADR/MAINSADR/n8691 ), .A(
        \SADR/MAINSADR/addindoff[15] ), .B(\SADR/m_fadrl[19] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U278  ( .ZN(\SADR/MAINSADR/n8831 ), .A(
        \SADR/pgaddwz[6] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[6] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[6] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[6] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_invx05 \SADR/MAINSADR/U344  ( .ZN(\SADR/MAINSADR/n8666 ), .A(
        \SADR/MAINSADR/n8662 ) );
    snl_invx05 \SADR/MAINSADR/U363  ( .ZN(\SADR/intbitno[3] ), .A(
        \SADR/MAINSADR/n8654 ) );
    snl_invx05 \SADR/MAINSADR/U101  ( .ZN(\SADR/MAINSADR/n8701 ), .A(
        \SADR/operand[25] ) );
    snl_muxi21x1 \SADR/MAINSADR/U231  ( .ZN(\SADR/MAINSADR/index[14] ), .A(
        \SADR/MAINSADR/n8892 ), .B(\SADR/MAINSADR/n8897 ), .S(ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U420  ( .ZN(\SADR/MAINSADR/oddadd[0] ), .A(
        \SADR/MAINSADR/n8664 ) );
    snl_nand04x0 \SADR/MAINSADR/U126  ( .ZN(\SADR/MAINSADR/n8730 ), .A(
        \SADR/MAINSADR/n8731 ), .B(\SADR/MAINSADR/n8732 ), .C(
        \SADR/MAINSADR/n8733 ), .D(\SADR/MAINSADR/n8734 ) );
    snl_and04x1 \SADR/MAINSADR/U211  ( .Z(\SADR/MAINSADR/n8854 ), .A(
        \SADR/MAINSADR/n8855 ), .B(\SADR/MAINSADR/n8856 ), .C(
        \SADR/MAINSADR/n8857 ), .D(\SADR/MAINSADR/n8858 ) );
    snl_and04x1 \SADR/MAINSADR/U216  ( .Z(\SADR/MAINSADR/n8863 ), .A(
        \SADR/MAINSADR/n8864 ), .B(\SADR/MAINSADR/n8865 ), .C(
        \SADR/MAINSADR/n8866 ), .D(\SADR/MAINSADR/n8867 ) );
    snl_nand02x1 \SADR/MAINSADR/U381  ( .ZN(\SADR/MAINSADR/n8770 ), .A(
        \SADR/MAINSADR/oddadd_p1[1] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_nand02x1 \SADR/MAINSADR/U386  ( .ZN(\SADR/MAINSADR/n8789 ), .A(
        \SADR/MAINSADR/oddadd_p1[14] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U407  ( .ZN(\SADR/MAINSADR/oddadd[6] ), .A(
        \SADR/MAINSADR/n8680 ) );
    snl_invx05 \SADR/MAINSADR/U400  ( .ZN(\SADR/MAINSADR/oddadd[12] ), .A(
        \SADR/MAINSADR/n8677 ) );
    snl_aoib122x0 \SADR/MAINSADR/U66  ( .ZN(\SADR/MAINSADR/n8671 ), .A(
        \SADR/MAINSADR/n8666 ), .B(\SADR/MAINSADR/oddadd[21] ), .C(
        \SADR/MAINSADR/oddadd_p1[21] ), .D(\SADR/MAINSADR/n8667 ), .E(
        \SADR/MAINSADR/n8672 ) );
    snl_and02x1 \SADR/MAINSADR/U106  ( .Z(\SADR/MAINSADR/n8706 ), .A(
        \SADR/MAINSADR/n8705 ), .B(\SADR/MAINSADR/n8702 ) );
    snl_and02x1 \SADR/MAINSADR/U121  ( .Z(\SADR/MAINSADR/n8721 ), .A(
        \SADR/MAINSADR/n8713 ), .B(\SADR/MAINSADR/n8709 ) );
    snl_and04x1 \SADR/MAINSADR/U236  ( .Z(\SADR/MAINSADR/n8912 ), .A(
        \SADR/MAINSADR/n8913 ), .B(\SADR/MAINSADR/n8914 ), .C(
        \SADR/MAINSADR/n8915 ), .D(\SADR/MAINSADR/n8916 ) );
    snl_invx05 \SADR/MAINSADR/U427  ( .ZN(\SADR/MAINSADR/oddadd[16] ), .A(
        \SADR/MAINSADR/n8690 ) );
    snl_muxi21x1 \SADR/MAINSADR/U83  ( .ZN(\SADR/MAINSADR/n8690 ), .A(
        \SADR/MAINSADR/addindoff[16] ), .B(\SADR/m_fadrl[20] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_muxi21x1 \SADR/MAINSADR/U168  ( .ZN(\pgregadrh[15] ), .A(
        \SADR/MAINSADR/n8797 ), .B(\SADR/MAINSADR/n8785 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi222x0 \SADR/MAINSADR/U258  ( .ZN(\SADR/MAINSADR/n8657 ), .A(
        \SADR/pgovfwxyz ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/MAINSADR/n8923 
        ), .D(\SADR/MAINSADR/n8643 ), .E(\SADR/sadr[27] ), .F(
        \SADR/MAINSADR/n8924 ) );
    snl_aoi222x0 \SADR/MAINSADR/U343  ( .ZN(\SADR/MAINSADR/n8913 ), .A(
        \pk_indw_h[10] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[10] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[10] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_nand02x1 \SADR/MAINSADR/U358  ( .ZN(\SADR/MAINSADR/n8650 ), .A(
        \SADR/MAINSADR/n8635 ), .B(\SADR/MAINSADR/oddadd[1] ) );
    snl_nor02x1 \SADR/MAINSADR/U364  ( .ZN(pgoddflgh), .A(
        \SADR/MAINSADR/n8695 ), .B(\SADR/MAINSADR/n8694 ) );
    snl_aoi222x0 \SADR/MAINSADR/U26  ( .ZN(\SADR/MAINSADR/n8799 ), .A(
        \SADR/MAINSADR/oddadd_m1[11] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[10] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[10] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U34  ( .ZN(\SADR/MAINSADR/n8771 ), .A(
        \SADR/MAINSADR/oddadd_m1[1] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[0] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[0] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_nand03x0 \SADR/MAINSADR/U98  ( .ZN(\SADR/MAINSADR/n8661 ), .A(
        \SADR/MAINSADR/n8696 ), .B(ph_lwdsrc_h), .C(ph_adrinc_h) );
    snl_oa112x1 \SADR/MAINSADR/U154  ( .Z(\SADR/MAINSADR/n8779 ), .A(
        \SADR/MAINSADR/n8689 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8780 ), .D(\SADR/MAINSADR/n8781 ) );
    snl_nor02x1 \SADR/MAINSADR/U48  ( .ZN(\SADR/MAINSADR/index[0] ), .A(
        ph_lwdsrc_h), .B(\SADR/MAINSADR/n8636 ) );
    snl_nand04x0 \SADR/MAINSADR/U128  ( .ZN(\SADR/MAINSADR/n8740 ), .A(
        \SADR/MAINSADR/n8741 ), .B(\SADR/MAINSADR/n8742 ), .C(
        \SADR/MAINSADR/n8743 ), .D(\SADR/MAINSADR/n8744 ) );
    snl_muxi21x1 \SADR/MAINSADR/U173  ( .ZN(\pgregadrh[11] ), .A(
        \SADR/MAINSADR/n8757 ), .B(\SADR/MAINSADR/n8797 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U243  ( .ZN(\SADR/MAINSADR/n8726 ), .A(
        \pk_indw_h[23] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[23] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[23] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U264  ( .ZN(\SADR/MAINSADR/n8818 ), .A(
        \SADR/pgaddwxyz[9] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[9] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[9] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[9] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_muxi21x1 \SADR/MAINSADR/U184  ( .ZN(\SADR/MAINSADR/offset[1] ), .A(
        \SADR/MAINSADR/n8809 ), .B(\SADR/MAINSADR/n8649 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_and04x1 \SADR/MAINSADR/U196  ( .Z(\SADR/MAINSADR/n8814 ), .A(
        \SADR/MAINSADR/n8815 ), .B(\SADR/MAINSADR/n8816 ), .C(
        \SADR/MAINSADR/n8817 ), .D(\SADR/MAINSADR/n8818 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U336  ( .ZN(\SADR/MAINSADR/n8911 ), .A(
        \SADR/pgaddwxyz[11] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[11] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[11] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[11] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U281  ( .ZN(\SADR/MAINSADR/n8837 ), .A(
        \SADR/pgaddwxy[5] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[5] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[5] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[5] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi222x0 \SADR/MAINSADR/U311  ( .ZN(\SADR/MAINSADR/n8873 ), .A(
        \pk_indw_h[18] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[18] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[18] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U324  ( .ZN(\SADR/MAINSADR/n8896 ), .A(
        \SADR/pgaddwxyz[14] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[14] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[14] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[14] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U293  ( .ZN(\SADR/MAINSADR/n8852 ), .A(
        \SADR/pgaddwxy[2] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[2] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[2] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[2] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi222x0 \SADR/MAINSADR/U303  ( .ZN(\SADR/MAINSADR/n8864 ), .A(
        \pk_indw_h[19] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[19] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[19] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi122x0 \SADR/MAINSADR/U146  ( .ZN(\SADR/MAINSADR/n8772 ), .A(
        \SADR/MAINSADR/oddadd_m1[0] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_p1[0] ), .D(\SADR/MAINSADR/n8667 ), .E(
        \SADR/MAINSADR/n8660 ) );
    snl_and04x1 \SADR/MAINSADR/U218  ( .Z(\SADR/MAINSADR/n8636 ), .A(
        \SADR/MAINSADR/n8868 ), .B(\SADR/MAINSADR/n8869 ), .C(
        \SADR/MAINSADR/n8870 ), .D(\SADR/MAINSADR/n8871 ) );
    snl_nand02x1 \SADR/MAINSADR/U388  ( .ZN(\SADR/MAINSADR/n8795 ), .A(
        \SADR/MAINSADR/oddadd_p1[12] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U409  ( .ZN(\SADR/MAINSADR/oddadd[9] ), .A(
        \SADR/MAINSADR/n8683 ) );
    snl_invx05 \SADR/MAINSADR/U91  ( .ZN(\SADR/MAINSADR/n8651 ), .A(
        \SADR/operand[2] ) );
    snl_oa112x1 \SADR/MAINSADR/U161  ( .Z(\SADR/MAINSADR/n8788 ), .A(
        \SADR/MAINSADR/n8692 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8789 ), .D(\SADR/MAINSADR/n8790 ) );
    snl_aoi222x0 \SADR/MAINSADR/U251  ( .ZN(\SADR/MAINSADR/n8736 ), .A(
        \pk_indw_h[21] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[21] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[21] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U276  ( .ZN(\SADR/MAINSADR/n8833 ), .A(
        \SADR/pgaddwxyz[6] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[6] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[6] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[6] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_and04x1 \SADR/MAINSADR/U203  ( .Z(\SADR/MAINSADR/n8834 ), .A(
        \SADR/MAINSADR/n8835 ), .B(\SADR/MAINSADR/n8836 ), .C(
        \SADR/MAINSADR/n8837 ), .D(\SADR/MAINSADR/n8838 ) );
    snl_invx05 \SADR/MAINSADR/U351  ( .ZN(\SADR/MAINSADR/n8803 ), .A(
        \SADR/operand[13] ) );
    snl_nand02x1 \SADR/MAINSADR/U376  ( .ZN(\SADR/MAINSADR/n8752 ), .A(
        \SADR/MAINSADR/oddadd_p1[8] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U393  ( .ZN(\SADR/MAINSADR/n8860 ), .A(
        \SADR/MAINSADR/n8730 ) );
    snl_invx05 \SADR/MAINSADR/U412  ( .ZN(\SADR/MAINSADR/oddadd[4] ), .A(
        \SADR/MAINSADR/n8684 ) );
    snl_aoi222x0 \SADR/MAINSADR/U20  ( .ZN(\SADR/MAINSADR/n8781 ), .A(
        \SADR/MAINSADR/oddadd_m1[17] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[16] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[16] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U27  ( .ZN(\SADR/MAINSADR/n8802 ), .A(
        \SADR/MAINSADR/oddadd_m1[10] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[9] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[9] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U35  ( .ZN(\SADR/MAINSADR/n8756 ), .A(
        \SADR/MAINSADR/oddadd_m1[4] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[3] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[3] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_ao012x1 \SADR/MAINSADR/U53  ( .Z(\SADR/MAINSADR/oddadd[23] ), .A(
        \SADR/MAINSADR/addindoff[23] ), .B(\SADR/MAINSADR/n8638 ), .C(
        \SADR/MAINSADR/n8639 ) );
    snl_muxi21x1 \SADR/MAINSADR/U74  ( .ZN(\SADR/MAINSADR/n8682 ), .A(
        \SADR/MAINSADR/addindoff[5] ), .B(\SADR/m_fadrl[9] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U114  ( .Z(\SADR/MAINSADR/n8714 ), .A(
        \SADR/MAINSADR/n8713 ), .B(\SADR/MAINSADR/n8702 ) );
    snl_oa112x1 \SADR/MAINSADR/U133  ( .Z(\SADR/MAINSADR/n8748 ), .A(
        \SADR/MAINSADR/n8682 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8749 ), .D(\SADR/MAINSADR/n8750 ) );
    snl_and04x1 \SADR/MAINSADR/U224  ( .Z(\SADR/MAINSADR/n8882 ), .A(
        \SADR/MAINSADR/n8883 ), .B(\SADR/MAINSADR/n8884 ), .C(
        \SADR/MAINSADR/n8885 ), .D(\SADR/MAINSADR/n8886 ) );
    snl_muxi21x1 \SADR/MAINSADR/U435  ( .ZN(\pgsdprlh[14] ), .A(
        \SADR/MAINSADR/n8681 ), .B(\SADR/MAINSADR/n8692 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_and02x1 \SADR/MAINSADR/U99  ( .Z(\SADR/MAINSADR/n8698 ), .A(
        ph_adrdec_h), .B(\SADR/MAINSADR/n8694 ) );
    snl_and04x1 \SADR/MAINSADR/U197  ( .Z(\SADR/MAINSADR/n8819 ), .A(
        \SADR/MAINSADR/n8820 ), .B(\SADR/MAINSADR/n8821 ), .C(
        \SADR/MAINSADR/n8822 ), .D(\SADR/MAINSADR/n8823 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U288  ( .ZN(\SADR/MAINSADR/n8848 ), .A(
        \SADR/pgaddwxyz[3] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[3] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[3] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[3] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U318  ( .ZN(\SADR/MAINSADR/n8884 ), .A(
        \SADR/pgaddwz[16] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[16] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[16] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[16] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U337  ( .ZN(\SADR/MAINSADR/n8910 ), .A(
        \SADR/pgaddwxy[11] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[11] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[11] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[11] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U280  ( .ZN(\SADR/MAINSADR/n8838 ), .A(
        \SADR/pgaddwxyz[5] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[5] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[5] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[5] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U310  ( .ZN(\SADR/MAINSADR/n8874 ), .A(
        \SADR/pgaddwz[18] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[18] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[18] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[18] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U155  ( .ZN(\pgregadrh[21] ), .A(
        \SADR/MAINSADR/n8779 ), .B(\SADR/MAINSADR/n8671 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_invx05 \SADR/MAINSADR/U359  ( .ZN(\SADR/intbitno[1] ), .A(
        \SADR/MAINSADR/n8650 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U265  ( .ZN(\SADR/MAINSADR/n8817 ), .A(
        \SADR/pgaddwxy[9] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[9] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[9] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[9] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_muxi21x2 \SADR/MAINSADR/U40  ( .ZN(\pgsdprlh[19] ), .A(
        \SADR/MAINSADR/n8691 ), .B(\SADR/MAINSADR/n8637 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U82  ( .ZN(\SADR/MAINSADR/n8689 ), .A(
        \SADR/MAINSADR/addindoff[17] ), .B(\SADR/m_fadrl[21] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_oa112x1 \SADR/MAINSADR/U169  ( .Z(\SADR/MAINSADR/n8800 ), .A(
        \SADR/MAINSADR/n8681 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8801 ), .D(\SADR/MAINSADR/n8802 ) );
    snl_muxi21x1 \SADR/MAINSADR/U172  ( .ZN(\pgregadrh[12] ), .A(
        \SADR/MAINSADR/n8751 ), .B(\SADR/MAINSADR/n8794 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U242  ( .ZN(\SADR/MAINSADR/n8727 ), .A(
        \SADR/pgaddwz[23] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[23] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[23] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[23] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi022x1 \SADR/MAINSADR/U259  ( .ZN(\SADR/MAINSADR/n8658 ), .A(
        \SADR/pgovfxyz ), .B(\SADR/MAINSADR/n8706 ), .C(\SADR/pgovfwyz ), .D(
        \SADR/MAINSADR/n8708 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U342  ( .ZN(\SADR/MAINSADR/n8914 ), .A(
        \SADR/pgaddwz[10] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[10] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[10] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[10] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_invx05 \SADR/MAINSADR/U365  ( .ZN(\SADR/MAINSADR/n8924 ), .A(
        \SADR/segbase[17] ) );
    snl_aoi012x1 \SADR/MAINSADR/U52  ( .ZN(\SADR/MAINSADR/n8642 ), .A(
        \SADR/MAINSADR/addindoff[22] ), .B(\SADR/MAINSADR/n8638 ), .C(
        \SADR/MAINSADR/n8639 ) );
    snl_aoib122x0 \SADR/MAINSADR/U67  ( .ZN(\SADR/MAINSADR/n8673 ), .A(
        \SADR/MAINSADR/n8666 ), .B(\SADR/MAINSADR/oddadd[20] ), .C(
        \SADR/MAINSADR/oddadd_p1[20] ), .D(\SADR/MAINSADR/n8667 ), .E(
        \SADR/MAINSADR/n8674 ) );
    snl_nor02x1 \SADR/MAINSADR/U107  ( .ZN(\SADR/MAINSADR/n8707 ), .A(
        \SADR/MAINSADR/n8700 ), .B(\SADR/operand[26] ) );
    snl_and02x1 \SADR/MAINSADR/U120  ( .Z(\SADR/MAINSADR/n8720 ), .A(
        \SADR/MAINSADR/n8719 ), .B(\SADR/MAINSADR/n8703 ) );
    snl_muxi21x1 \SADR/MAINSADR/U210  ( .ZN(\SADR/MAINSADR/index[3] ), .A(
        \SADR/MAINSADR/n8844 ), .B(\SADR/MAINSADR/n8849 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U380  ( .ZN(\SADR/MAINSADR/n8764 ), .A(
        \SADR/MAINSADR/oddadd_p1[6] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U401  ( .ZN(\SADR/MAINSADR/oddadd[8] ), .A(
        \SADR/MAINSADR/n8675 ) );
    snl_muxi21x1 \SADR/MAINSADR/U237  ( .ZN(\SADR/MAINSADR/index[11] ), .A(
        \SADR/MAINSADR/n8907 ), .B(\SADR/MAINSADR/n8912 ), .S(ph_lwdsrc_h) );
    snl_muxi21x1 \SADR/MAINSADR/U426  ( .ZN(\pgsdprlh[21] ), .A(
        \SADR/MAINSADR/n8689 ), .B(\SADR/MAINSADR/n8641 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U75  ( .ZN(\SADR/MAINSADR/n8683 ), .A(
        \SADR/MAINSADR/addindoff[9] ), .B(\SADR/m_fadrl[13] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U115  ( .Z(\SADR/MAINSADR/n8715 ), .A(
        \SADR/MAINSADR/n8709 ), .B(\SADR/MAINSADR/n8705 ) );
    snl_oa112x1 \SADR/MAINSADR/U132  ( .Z(\SADR/MAINSADR/n8745 ), .A(
        \SADR/MAINSADR/n8683 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8746 ), .D(\SADR/MAINSADR/n8747 ) );
    snl_muxi21x1 \SADR/MAINSADR/U202  ( .ZN(\SADR/MAINSADR/index[7] ), .A(
        \SADR/MAINSADR/n8824 ), .B(\SADR/MAINSADR/n8829 ), .S(ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U392  ( .ZN(\SADR/MAINSADR/n8861 ), .A(
        \SADR/MAINSADR/n8735 ) );
    snl_muxi21x1 \SADR/MAINSADR/U413  ( .ZN(\pgsdprlh[8] ), .A(
        \SADR/MAINSADR/n8684 ), .B(\SADR/MAINSADR/n8675 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_invx05 \SADR/MAINSADR/U90  ( .ZN(\SADR/MAINSADR/n8653 ), .A(
        \SADR/operand[3] ) );
    snl_muxi21x1 \SADR/MAINSADR/U225  ( .ZN(\SADR/MAINSADR/index[17] ), .A(
        \SADR/MAINSADR/n8877 ), .B(\SADR/MAINSADR/n8882 ), .S(ph_lwdsrc_h) );
    snl_aoi2222x0 \SADR/MAINSADR/U289  ( .ZN(\SADR/MAINSADR/n8847 ), .A(
        \SADR/pgaddwxy[3] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[3] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[3] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[3] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi222x0 \SADR/MAINSADR/U319  ( .ZN(\SADR/MAINSADR/n8883 ), .A(
        \pk_indw_h[16] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[16] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[16] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U434  ( .ZN(\pgsdprlh[16] ), .A(
        \SADR/MAINSADR/n8677 ), .B(\SADR/MAINSADR/n8690 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_invx05 \SADR/MAINSADR/U350  ( .ZN(\SADR/MAINSADR/n8805 ), .A(
        \SADR/operand[12] ) );
    snl_muxi21x1 \SADR/MAINSADR/U147  ( .ZN(\pgregadrh[4] ), .A(
        \SADR/MAINSADR/n8772 ), .B(\SADR/MAINSADR/n8754 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_nand02x1 \SADR/MAINSADR/U377  ( .ZN(\SADR/MAINSADR/n8761 ), .A(
        \SADR/MAINSADR/oddadd_p1[3] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U277  ( .ZN(\SADR/MAINSADR/n8832 ), .A(
        \SADR/pgaddwxy[6] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[6] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[6] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[6] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi012x1 \SADR/MAINSADR/U49  ( .ZN(\SADR/MAINSADR/n8637 ), .A(
        \SADR/MAINSADR/addindoff[19] ), .B(\SADR/MAINSADR/n8638 ), .C(
        \SADR/MAINSADR/n8639 ) );
    snl_invx05 \SADR/MAINSADR/U129  ( .ZN(\SADR/MAINSADR/n8646 ), .A(
        \SADR/operand[22] ) );
    snl_muxi21x1 \SADR/MAINSADR/U160  ( .ZN(\pgregadrh[19] ), .A(
        \SADR/MAINSADR/n8785 ), .B(\SADR/MAINSADR/n8773 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U250  ( .ZN(\SADR/MAINSADR/n8737 ), .A(
        \SADR/pgaddwz[21] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[21] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[21] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[21] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_mux21x1 \SADR/MAINSADR/U185  ( .Z(\SADR/MAINSADR/offset[19] ), .A(
        \SADR/operand[23] ), .B(\SADR/operand[19] ), .S(\SADR/MAINSADR/n8634 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U325  ( .ZN(\SADR/MAINSADR/n8895 ), .A(
        \SADR/pgaddwxy[14] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[14] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[14] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[14] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U292  ( .ZN(\SADR/MAINSADR/n8853 ), .A(
        \SADR/pgaddwxyz[2] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[2] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[2] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[2] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U302  ( .ZN(\SADR/MAINSADR/n8865 ), .A(
        \SADR/pgaddwz[19] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[19] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[19] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[19] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U219  ( .ZN(\SADR/MAINSADR/index[1] ), .A(
        \SADR/MAINSADR/n8854 ), .B(\SADR/MAINSADR/n8636 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U389  ( .ZN(\SADR/MAINSADR/n8798 ), .A(
        \SADR/MAINSADR/oddadd_p1[11] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_muxi21x1 \SADR/MAINSADR/U408  ( .ZN(\pgsdprlh[10] ), .A(
        \SADR/MAINSADR/n8680 ), .B(\SADR/MAINSADR/n8681 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U69  ( .ZN(\SADR/MAINSADR/n8677 ), .A(
        \SADR/MAINSADR/addindoff[12] ), .B(\SADR/m_fadrl[16] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U109  ( .Z(\SADR/MAINSADR/n8709 ), .A(
        \SADR/operand[24] ), .B(\SADR/MAINSADR/n8701 ) );
    snl_mux21x1 \SADR/MAINSADR/U182  ( .Z(\SADR/MAINSADR/offset[3] ), .A(
        \SADR/operand[7] ), .B(\SADR/operand[3] ), .S(\SADR/MAINSADR/n8634 )
         );
    snl_aoi222x0 \SADR/MAINSADR/U295  ( .ZN(\SADR/MAINSADR/n8850 ), .A(
        \pk_indw_h[2] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[2] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[2] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U305  ( .ZN(\SADR/MAINSADR/n8870 ), .A(
        \SADR/pgaddwxy[0] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[0] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[0] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[0] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U322  ( .ZN(\SADR/MAINSADR/n8889 ), .A(
        \SADR/pgaddwz[15] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[15] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[15] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[15] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_oa112x1 \SADR/MAINSADR/U167  ( .Z(\SADR/MAINSADR/n8797 ), .A(
        \SADR/MAINSADR/n8679 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8798 ), .D(\SADR/MAINSADR/n8799 ) );
    snl_aoi022x1 \SADR/MAINSADR/U239  ( .ZN(\SADR/MAINSADR/n8774 ), .A(
        \SADR/MAINSADR/oddadd_p1[19] ), .B(\SADR/MAINSADR/n8667 ), .C(
        \SADR/MAINSADR/n8666 ), .D(\SADR/MAINSADR/oddadd[19] ) );
    snl_muxi21x1 \SADR/MAINSADR/U428  ( .ZN(\pgsdprlh[20] ), .A(
        \SADR/MAINSADR/n8690 ), .B(\SADR/MAINSADR/n8640 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_oai113x0 \SADR/MAINSADR/U257  ( .ZN(\SADR/MAINSADR/n8656 ), .A(
        \SADR/MAINSADR/n8694 ), .B(\SADR/MAINSADR/n8920 ), .C(
        \SADR/MAINSADR/n8921 ), .D(\SADR/MAINSADR/n8922 ), .E(
        \SADR/MAINSADR/n8919 ) );
    snl_aoi222x0 \SADR/MAINSADR/U29  ( .ZN(\SADR/MAINSADR/n8753 ), .A(
        \SADR/MAINSADR/oddadd_m1[8] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[7] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[7] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_nand14x2 \SADR/MAINSADR/U47  ( .ZN(pgadrovfh), .A(
        \SADR/MAINSADR/n8656 ), .B(\SADR/MAINSADR/n8657 ), .C(
        \SADR/MAINSADR/n8658 ), .D(\SADR/MAINSADR/n8659 ) );
    snl_nor02x1 \SADR/MAINSADR/U55  ( .ZN(\SADR/MAINSADR/offset[21] ), .A(
        \SADR/MAINSADR/n8643 ), .B(\SADR/MAINSADR/n8645 ) );
    snl_muxi21x1 \SADR/MAINSADR/U72  ( .ZN(\SADR/MAINSADR/n8680 ), .A(
        \SADR/MAINSADR/addindoff[6] ), .B(\SADR/m_fadrl[10] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_invx05 \SADR/MAINSADR/U97  ( .ZN(\SADR/MAINSADR/n8697 ), .A(
        ph_adrinc_h) );
    snl_muxi21x1 \SADR/MAINSADR/U140  ( .ZN(\pgregadrh[7] ), .A(
        \SADR/MAINSADR/n8760 ), .B(\SADR/MAINSADR/n8757 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U270  ( .ZN(\SADR/MAINSADR/n8821 ), .A(
        \SADR/pgaddwz[8] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[8] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[8] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[8] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_invx05 \SADR/MAINSADR/U370  ( .ZN(\SADR/MAINSADR/oddadd[21] ), .A(
        \SADR/MAINSADR/n8641 ) );
    snl_and04x1 \SADR/MAINSADR/U222  ( .Z(\SADR/MAINSADR/n8877 ), .A(
        \SADR/MAINSADR/n8878 ), .B(\SADR/MAINSADR/n8879 ), .C(
        \SADR/MAINSADR/n8880 ), .D(\SADR/MAINSADR/n8881 ) );
    snl_invx05 \SADR/MAINSADR/U357  ( .ZN(\SADR/intbitno[0] ), .A(
        \SADR/MAINSADR/n8648 ) );
    snl_muxi21x1 \SADR/MAINSADR/U433  ( .ZN(\pgsdprlh[17] ), .A(
        \SADR/MAINSADR/n8693 ), .B(\SADR/MAINSADR/n8689 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_and02x1 \SADR/MAINSADR/U112  ( .Z(\SADR/MAINSADR/n8712 ), .A(
        \SADR/MAINSADR/n8711 ), .B(\SADR/MAINSADR/n8703 ) );
    snl_oa112x1 \SADR/MAINSADR/U135  ( .Z(\SADR/MAINSADR/n8751 ), .A(
        \SADR/MAINSADR/n8675 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8752 ), .D(\SADR/MAINSADR/n8753 ) );
    snl_and04x1 \SADR/MAINSADR/U205  ( .Z(\SADR/MAINSADR/n8839 ), .A(
        \SADR/MAINSADR/n8840 ), .B(\SADR/MAINSADR/n8841 ), .C(
        \SADR/MAINSADR/n8842 ), .D(\SADR/MAINSADR/n8843 ) );
    snl_nor04x0 \SADR/MAINSADR/U395  ( .ZN(\SADR/MAINSADR/n8920 ), .A(
        \SADR/MAINSADR/n8740 ), .B(\SADR/MAINSADR/n8735 ), .C(
        \SADR/MAINSADR/n8730 ), .D(\SADR/MAINSADR/n8725 ) );
    snl_invx05 \SADR/MAINSADR/U414  ( .ZN(\SADR/MAINSADR/oddadd[3] ), .A(
        \SADR/MAINSADR/n8685 ) );
    snl_oai012x1 \SADR/MAINSADR/U60  ( .ZN(\pgsdprlh[2] ), .A(
        \SADR/MAINSADR/n8634 ), .B(\SADR/MAINSADR/n8651 ), .C(
        \SADR/MAINSADR/n8652 ) );
    snl_and04x1 \SADR/MAINSADR/U199  ( .Z(\SADR/MAINSADR/n8824 ), .A(
        \SADR/MAINSADR/n8825 ), .B(\SADR/MAINSADR/n8826 ), .C(
        \SADR/MAINSADR/n8827 ), .D(\SADR/MAINSADR/n8828 ) );
    snl_aoi222x0 \SADR/MAINSADR/U339  ( .ZN(\SADR/MAINSADR/n8908 ), .A(
        \pk_indw_h[11] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[11] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[11] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_and04x1 \SADR/MAINSADR/U230  ( .Z(\SADR/MAINSADR/n8897 ), .A(
        \SADR/MAINSADR/n8898 ), .B(\SADR/MAINSADR/n8899 ), .C(
        \SADR/MAINSADR/n8900 ), .D(\SADR/MAINSADR/n8901 ) );
    snl_muxi21x1 \SADR/MAINSADR/U421  ( .ZN(\pgsdprlh[4] ), .A(
        \SADR/MAINSADR/n8664 ), .B(\SADR/MAINSADR/n8684 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_invx05 \SADR/MAINSADR/U100  ( .ZN(\SADR/MAINSADR/n8700 ), .A(
        \SADR/operand[27] ) );
    snl_nand04x0 \SADR/MAINSADR/U127  ( .ZN(\SADR/MAINSADR/n8735 ), .A(
        \SADR/MAINSADR/n8736 ), .B(\SADR/MAINSADR/n8737 ), .C(
        \SADR/MAINSADR/n8738 ), .D(\SADR/MAINSADR/n8739 ) );
    snl_muxi21x1 \SADR/MAINSADR/U217  ( .ZN(\SADR/MAINSADR/index[20] ), .A(
        \SADR/MAINSADR/n8862 ), .B(\SADR/MAINSADR/n8863 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U387  ( .ZN(\SADR/MAINSADR/n8792 ), .A(
        \SADR/MAINSADR/oddadd_p1[13] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U406  ( .ZN(\SADR/MAINSADR/oddadd[10] ), .A(
        \SADR/MAINSADR/n8681 ) );
    snl_muxi21x1 \SADR/MAINSADR/U149  ( .ZN(\pgregadrh[2] ), .A(
        \SADR/MAINSADR/n8651 ), .B(\SADR/MAINSADR/n8766 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U279  ( .ZN(\SADR/MAINSADR/n8830 ), .A(
        \pk_indw_h[6] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[6] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[6] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U85  ( .ZN(\SADR/MAINSADR/n8692 ), .A(
        \SADR/MAINSADR/addindoff[14] ), .B(\SADR/m_fadrl[18] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_nand02x1 \SADR/MAINSADR/U362  ( .ZN(\SADR/MAINSADR/n8654 ), .A(
        \SADR/MAINSADR/n8635 ), .B(\SADR/MAINSADR/oddadd[3] ) );
    snl_invx05 \SADR/MAINSADR/U345  ( .ZN(\SADR/MAINSADR/n8809 ), .A(
        \SADR/operand[5] ) );
    snl_nand02x1 \SADR/MAINSADR/U379  ( .ZN(\SADR/MAINSADR/n8767 ), .A(
        \SADR/MAINSADR/oddadd_p1[2] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_aoi222x0 \SADR/MAINSADR/U15  ( .ZN(\SADR/MAINSADR/n8670 ), .A(
        \SADR/MAINSADR/oddadd_m1[22] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[21] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[21] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_muxi21x1 \SADR/MAINSADR/U175  ( .ZN(\pgregadrh[0] ), .A(
        \SADR/MAINSADR/n8647 ), .B(\SADR/MAINSADR/n8772 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U17  ( .ZN(\SADR/MAINSADR/n8674 ), .A(
        \SADR/MAINSADR/oddadd_m1[20] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[19] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[19] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U22  ( .ZN(\SADR/MAINSADR/n8787 ), .A(
        \SADR/MAINSADR/oddadd_m1[15] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[14] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[14] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U32  ( .ZN(\SADR/MAINSADR/n8768 ), .A(
        \SADR/MAINSADR/oddadd_m1[2] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[1] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[1] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U245  ( .ZN(\SADR/MAINSADR/n8733 ), .A(
        \SADR/pgaddwxy[22] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[22] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[22] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[22] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_invx2 \SADR/MAINSADR/U39  ( .ZN(\SADR/MAINSADR/n8635 ), .A(
        \SADR/MAINSADR/n8633 ) );
    snl_and02x1 \SADR/MAINSADR/U57  ( .Z(\SADR/MAINSADR/offset[23] ), .A(
        \SADR/MAINSADR/n8635 ), .B(\SADR/operand[23] ) );
    snl_muxi21x1 \SADR/MAINSADR/U137  ( .ZN(\pgregadrh[8] ), .A(
        \SADR/MAINSADR/n8754 ), .B(\SADR/MAINSADR/n8751 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_oa112x1 \SADR/MAINSADR/U152  ( .Z(\SADR/MAINSADR/n8776 ), .A(
        \SADR/MAINSADR/n8688 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8777 ), .D(\SADR/MAINSADR/n8778 ) );
    snl_aoi022x1 \SADR/MAINSADR/U262  ( .ZN(\SADR/MAINSADR/n8927 ), .A(
        \SADR/pgovfwz ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgovfwy ), .D(
        \SADR/MAINSADR/n8718 ) );
    snl_muxi21x1 \SADR/MAINSADR/U190  ( .ZN(\SADR/MAINSADR/offset[14] ), .A(
        \SADR/MAINSADR/n8810 ), .B(\SADR/MAINSADR/n8813 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U287  ( .ZN(\SADR/MAINSADR/n8840 ), .A(
        \pk_indw_h[4] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[4] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[4] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U317  ( .ZN(\SADR/MAINSADR/n8885 ), .A(
        \SADR/pgaddwxy[16] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[16] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[16] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[16] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U330  ( .ZN(\SADR/MAINSADR/n8899 ), .A(
        \SADR/pgaddwz[13] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[13] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[13] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[13] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U70  ( .ZN(\SADR/MAINSADR/n8678 ), .A(
        \SADR/MAINSADR/addindoff[7] ), .B(\SADR/m_fadrl[11] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and04x1 \SADR/MAINSADR/U207  ( .Z(\SADR/MAINSADR/n8844 ), .A(
        \SADR/MAINSADR/n8845 ), .B(\SADR/MAINSADR/n8846 ), .C(
        \SADR/MAINSADR/n8847 ), .D(\SADR/MAINSADR/n8848 ) );
    snl_nor04x0 \SADR/MAINSADR/U397  ( .ZN(\SADR/MAINSADR/n8921 ), .A(
        \SADR/MAINSADR/n8859 ), .B(\SADR/MAINSADR/n8860 ), .C(
        \SADR/MAINSADR/n8861 ), .D(\SADR/MAINSADR/n8862 ) );
    snl_invx05 \SADR/MAINSADR/U416  ( .ZN(\SADR/MAINSADR/oddadd[2] ), .A(
        \SADR/MAINSADR/n8686 ) );
    snl_and02x1 \SADR/MAINSADR/U110  ( .Z(\SADR/MAINSADR/n8710 ), .A(
        \SADR/MAINSADR/n8709 ), .B(\SADR/MAINSADR/n8703 ) );
    snl_and04x1 \SADR/MAINSADR/U220  ( .Z(\SADR/MAINSADR/n8872 ), .A(
        \SADR/MAINSADR/n8873 ), .B(\SADR/MAINSADR/n8874 ), .C(
        \SADR/MAINSADR/n8875 ), .D(\SADR/MAINSADR/n8876 ) );
    snl_muxi21x1 \SADR/MAINSADR/U431  ( .ZN(\pgsdprlh[18] ), .A(
        \SADR/MAINSADR/n8692 ), .B(\SADR/MAINSADR/n8688 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_oa112x1 \SADR/MAINSADR/U159  ( .Z(\SADR/MAINSADR/n8785 ), .A(
        \SADR/MAINSADR/n8691 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8786 ), .D(\SADR/MAINSADR/n8787 ) );
    snl_nor02x1 \SADR/MAINSADR/U95  ( .ZN(\SADR/MAINSADR/n8696 ), .A(
        pgfbadrsel), .B(pgoddflgh) );
    snl_aoi2222x0 \SADR/MAINSADR/U269  ( .ZN(\SADR/MAINSADR/n8822 ), .A(
        \SADR/pgaddwxy[8] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[8] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[8] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[8] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_invx05 \SADR/MAINSADR/U355  ( .ZN(\SADR/MAINSADR/n8810 ), .A(
        \SADR/operand[18] ) );
    snl_aoi2222x0 \SADR/MAINSADR/U272  ( .ZN(\SADR/MAINSADR/n8828 ), .A(
        \SADR/pgaddwxyz[7] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[7] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[7] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[7] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_invx05 \SADR/MAINSADR/U369  ( .ZN(\SADR/MAINSADR/oddadd[22] ), .A(
        \SADR/MAINSADR/n8642 ) );
    snl_nand12x1 \SADR/MAINSADR/U372  ( .ZN(\SADR/MAINSADR/n8699 ), .A(
        \SADR/MAINSADR/n8696 ), .B(ph_lwdsrc_h) );
    snl_aoi222x0 \SADR/MAINSADR/U30  ( .ZN(\SADR/MAINSADR/n8759 ), .A(
        \SADR/MAINSADR/oddadd_m1[7] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[6] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[6] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_muxi21x1 \SADR/MAINSADR/U79  ( .ZN(\SADR/MAINSADR/n8687 ), .A(
        \SADR/MAINSADR/addindoff[1] ), .B(\SADR/m_fadrl[5] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_nor02x1 \SADR/MAINSADR/U119  ( .ZN(\SADR/MAINSADR/n8719 ), .A(
        \SADR/operand[24] ), .B(\SADR/operand[25] ) );
    snl_oa112x1 \SADR/MAINSADR/U142  ( .Z(\SADR/MAINSADR/n8766 ), .A(
        \SADR/MAINSADR/n8686 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8767 ), .D(\SADR/MAINSADR/n8768 ) );
    snl_oa112x1 \SADR/MAINSADR/U165  ( .Z(\SADR/MAINSADR/n8794 ), .A(
        \SADR/MAINSADR/n8677 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8795 ), .D(\SADR/MAINSADR/n8796 ) );
    snl_muxi21x1 \SADR/MAINSADR/U180  ( .ZN(\SADR/MAINSADR/offset[5] ), .A(
        \SADR/MAINSADR/n8804 ), .B(\SADR/MAINSADR/n8809 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi222x0 \SADR/MAINSADR/U255  ( .ZN(\SADR/MAINSADR/n8741 ), .A(
        \SADR/MAINSADR/n8724 ), .B(\pk_indw_h[20] ), .C(\SADR/MAINSADR/n8722 ), 
        .D(\pk_indy_h[20] ), .E(\SADR/MAINSADR/n8723 ), .F(\pk_indx_h[20] ) );
    snl_muxi21x1 \SADR/MAINSADR/U192  ( .ZN(\SADR/MAINSADR/offset[12] ), .A(
        \SADR/MAINSADR/n8812 ), .B(\SADR/MAINSADR/n8805 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U297  ( .ZN(\SADR/MAINSADR/n8857 ), .A(
        \SADR/pgaddwxy[1] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[1] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[1] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[1] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U320  ( .ZN(\SADR/MAINSADR/n8891 ), .A(
        \SADR/pgaddwxyz[15] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[15] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[15] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[15] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi222x0 \SADR/MAINSADR/U307  ( .ZN(\SADR/MAINSADR/n8868 ), .A(
        \pk_indw_h[0] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[0] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[0] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U285  ( .ZN(\SADR/MAINSADR/n8842 ), .A(
        \SADR/pgaddwxy[4] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[4] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[4] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[4] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi222x0 \SADR/MAINSADR/U315  ( .ZN(\SADR/MAINSADR/n8878 ), .A(
        \pk_indw_h[17] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[17] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[17] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U332  ( .ZN(\SADR/MAINSADR/n8906 ), .A(
        \SADR/pgaddwxyz[12] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[12] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[12] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[12] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_muxi21x1 \SADR/MAINSADR/U229  ( .ZN(\SADR/MAINSADR/index[15] ), .A(
        \SADR/MAINSADR/n8887 ), .B(\SADR/MAINSADR/n8892 ), .S(ph_lwdsrc_h) );
    snl_aoi222x0 \SADR/MAINSADR/U260  ( .ZN(\SADR/MAINSADR/n8925 ), .A(
        \SADR/pgovfyz ), .B(\SADR/MAINSADR/n8714 ), .C(\SADR/pgovfwxz ), .D(
        \SADR/MAINSADR/n8710 ), .E(\SADR/pgovfwxy ), .F(\SADR/MAINSADR/n8712 )
         );
    snl_and02x1 \SADR/MAINSADR/U150  ( .Z(\SADR/MAINSADR/n8773 ), .A(
        \SADR/MAINSADR/n8774 ), .B(\SADR/MAINSADR/n8775 ) );
    snl_muxi21x1 \SADR/MAINSADR/U177  ( .ZN(\SADR/MAINSADR/offset[8] ), .A(
        \SADR/MAINSADR/n8805 ), .B(\SADR/MAINSADR/n8806 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U247  ( .ZN(\SADR/MAINSADR/n8731 ), .A(
        \pk_indw_h[22] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[22] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[22] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi222x0 \SADR/MAINSADR/U45  ( .ZN(\SADR/MAINSADR/n8765 ), .A(
        \SADR/MAINSADR/oddadd_m1[6] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[5] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[5] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_invx05 \SADR/MAINSADR/U87  ( .ZN(\SADR/MAINSADR/n8655 ), .A(pgfbadrsel
        ) );
    snl_invx05 \SADR/MAINSADR/U347  ( .ZN(\SADR/MAINSADR/n8806 ), .A(
        \SADR/operand[8] ) );
    snl_nand04x0 \SADR/MAINSADR/U125  ( .ZN(\SADR/MAINSADR/n8725 ), .A(
        \SADR/MAINSADR/n8726 ), .B(\SADR/MAINSADR/n8727 ), .C(
        \SADR/MAINSADR/n8728 ), .D(\SADR/MAINSADR/n8729 ) );
    snl_nand02x1 \SADR/MAINSADR/U360  ( .ZN(\SADR/MAINSADR/n8652 ), .A(
        \SADR/MAINSADR/n8634 ), .B(\SADR/MAINSADR/oddadd[2] ) );
    snl_aoi222x0 \SADR/MAINSADR/U19  ( .ZN(\SADR/MAINSADR/n8778 ), .A(
        \SADR/MAINSADR/oddadd_m1[18] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[17] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[17] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U25  ( .ZN(\SADR/MAINSADR/n8796 ), .A(
        \SADR/MAINSADR/oddadd_m1[12] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[11] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[11] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_invx05 \SADR/MAINSADR/U37  ( .ZN(\SADR/MAINSADR/n8633 ), .A(
        ph_bitsrc_h) );
    snl_nand13x2 \SADR/MAINSADR/U42  ( .ZN(\SADR/MAINSADR/n8662 ), .A(
        ph_adrdec_h), .B(\SADR/MAINSADR/n8697 ), .C(\SADR/MAINSADR/n8699 ) );
    snl_oai012x1 \SADR/MAINSADR/U62  ( .ZN(\SADR/sadr[0] ), .A(ph_lwdsrc_h), 
        .B(\pgsdprlh[4] ), .C(\SADR/MAINSADR/n8655 ) );
    snl_muxi21x1 \SADR/MAINSADR/U215  ( .ZN(\SADR/MAINSADR/index[21] ), .A(
        \SADR/MAINSADR/n8861 ), .B(\SADR/MAINSADR/n8862 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U385  ( .ZN(\SADR/MAINSADR/n8786 ), .A(
        \SADR/MAINSADR/oddadd_p1[15] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U404  ( .ZN(\SADR/MAINSADR/oddadd[7] ), .A(
        \SADR/MAINSADR/n8678 ) );
    snl_aoib122x0 \SADR/MAINSADR/U65  ( .ZN(\SADR/MAINSADR/n8669 ), .A(
        \SADR/MAINSADR/n8666 ), .B(\SADR/MAINSADR/oddadd[22] ), .C(
        \SADR/MAINSADR/oddadd_p1[22] ), .D(\SADR/MAINSADR/n8667 ), .E(
        \SADR/MAINSADR/n8670 ) );
    snl_and02x1 \SADR/MAINSADR/U102  ( .Z(\SADR/MAINSADR/n8702 ), .A(
        \SADR/operand[25] ), .B(\SADR/operand[24] ) );
    snl_and04x1 \SADR/MAINSADR/U232  ( .Z(\SADR/MAINSADR/n8902 ), .A(
        \SADR/MAINSADR/n8903 ), .B(\SADR/MAINSADR/n8904 ), .C(
        \SADR/MAINSADR/n8905 ), .D(\SADR/MAINSADR/n8906 ) );
    snl_invx05 \SADR/MAINSADR/U423  ( .ZN(\SADR/MAINSADR/oddadd[18] ), .A(
        \SADR/MAINSADR/n8688 ) );
    snl_and02x1 \SADR/MAINSADR/U105  ( .Z(\SADR/MAINSADR/n8705 ), .A(
        \SADR/operand[26] ), .B(\SADR/MAINSADR/n8700 ) );
    snl_mux21x1 \SADR/MAINSADR/U189  ( .Z(\SADR/MAINSADR/offset[15] ), .A(
        \SADR/operand[19] ), .B(\SADR/operand[15] ), .S(\SADR/MAINSADR/n8634 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U329  ( .ZN(\SADR/MAINSADR/n8900 ), .A(
        \SADR/pgaddwxy[13] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[13] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[13] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[13] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_muxi21x1 \SADR/MAINSADR/U235  ( .ZN(\SADR/MAINSADR/index[12] ), .A(
        \SADR/MAINSADR/n8902 ), .B(\SADR/MAINSADR/n8907 ), .S(ph_lwdsrc_h) );
    snl_muxi21x1 \SADR/MAINSADR/U424  ( .ZN(\pgsdprlh[22] ), .A(
        \SADR/MAINSADR/n8688 ), .B(\SADR/MAINSADR/n8642 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U212  ( .ZN(\SADR/MAINSADR/index[2] ), .A(
        \SADR/MAINSADR/n8849 ), .B(\SADR/MAINSADR/n8854 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U382  ( .ZN(\SADR/MAINSADR/n8777 ), .A(
        \SADR/MAINSADR/oddadd_p1[18] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_invx05 \SADR/MAINSADR/U403  ( .ZN(\SADR/MAINSADR/oddadd[11] ), .A(
        \SADR/MAINSADR/n8679 ) );
    snl_muxi21x1 \SADR/MAINSADR/U80  ( .ZN(\SADR/MAINSADR/n8664 ), .A(
        \SADR/MAINSADR/addindoff[0] ), .B(\SADR/m_fadrl[4] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U122  ( .Z(\SADR/MAINSADR/n8722 ), .A(
        \SADR/MAINSADR/n8713 ), .B(\SADR/MAINSADR/n8711 ) );
    snl_aoi222x0 \SADR/MAINSADR/U299  ( .ZN(\SADR/MAINSADR/n8855 ), .A(
        \pk_indw_h[1] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[1] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[1] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U309  ( .ZN(\SADR/MAINSADR/n8875 ), .A(
        \SADR/pgaddwxy[18] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[18] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[18] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[18] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_invx05 \SADR/MAINSADR/U367  ( .ZN(\SADR/MAINSADR/n8638 ), .A(
        \SADR/MAINSADR/n8676 ) );
    snl_muxi21x1 \SADR/MAINSADR/U157  ( .ZN(\pgregadrh[20] ), .A(
        \SADR/MAINSADR/n8782 ), .B(\SADR/MAINSADR/n8673 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U170  ( .ZN(\pgregadrh[14] ), .A(
        \SADR/MAINSADR/n8800 ), .B(\SADR/MAINSADR/n8788 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U240  ( .ZN(\SADR/MAINSADR/n8729 ), .A(
        \SADR/pgaddwxyz[23] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[23] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[23] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[23] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U340  ( .ZN(\SADR/MAINSADR/n8916 ), .A(
        \SADR/pgaddwxyz[10] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[10] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[10] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[10] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_oai012x1 \SADR/MAINSADR/U59  ( .ZN(\pgsdprlh[1] ), .A(
        \SADR/MAINSADR/n8634 ), .B(\SADR/MAINSADR/n8649 ), .C(
        \SADR/MAINSADR/n8650 ) );
    snl_oa112x1 \SADR/MAINSADR/U139  ( .Z(\SADR/MAINSADR/n8760 ), .A(
        \SADR/MAINSADR/n8685 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8761 ), .D(\SADR/MAINSADR/n8762 ) );
    snl_muxi21x1 \SADR/MAINSADR/U195  ( .ZN(\SADR/MAINSADR/offset[0] ), .A(
        \SADR/MAINSADR/n8695 ), .B(\SADR/MAINSADR/n8647 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U267  ( .ZN(\SADR/MAINSADR/n8815 ), .A(
        \pk_indw_h[9] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[9] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[9] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U282  ( .ZN(\SADR/MAINSADR/n8836 ), .A(
        \SADR/pgaddwz[5] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[5] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[5] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[5] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U312  ( .ZN(\SADR/MAINSADR/n8881 ), .A(
        \SADR/pgaddwxyz[17] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[17] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[17] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[17] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_aoi222x0 \SADR/MAINSADR/U335  ( .ZN(\SADR/MAINSADR/n8903 ), .A(
        \pk_indw_h[12] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[12] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[12] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_invx05 \SADR/MAINSADR/U89  ( .ZN(\SADR/MAINSADR/n8643 ), .A(
        \SADR/MAINSADR/n8634 ) );
    snl_muxi21x1 \SADR/MAINSADR/U187  ( .ZN(\SADR/MAINSADR/offset[17] ), .A(
        \SADR/MAINSADR/n8645 ), .B(\SADR/MAINSADR/n8811 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_and04x1 \SADR/MAINSADR/U209  ( .Z(\SADR/MAINSADR/n8849 ), .A(
        \SADR/MAINSADR/n8850 ), .B(\SADR/MAINSADR/n8851 ), .C(
        \SADR/MAINSADR/n8852 ), .D(\SADR/MAINSADR/n8853 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U290  ( .ZN(\SADR/MAINSADR/n8846 ), .A(
        \SADR/pgaddwz[3] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[3] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[3] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[3] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U300  ( .ZN(\SADR/MAINSADR/n8867 ), .A(
        \SADR/pgaddwxyz[19] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[19] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[19] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[19] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_nand02x1 \SADR/MAINSADR/U399  ( .ZN(\SADR/MAINSADR/n8928 ), .A(
        \SADR/pgovfwx ), .B(\SADR/MAINSADR/n8720 ) );
    snl_invx05 \SADR/MAINSADR/U418  ( .ZN(\SADR/MAINSADR/oddadd[1] ), .A(
        \SADR/MAINSADR/n8687 ) );
    snl_aoi222x0 \SADR/MAINSADR/U327  ( .ZN(\SADR/MAINSADR/n8893 ), .A(
        \pk_indw_h[14] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[14] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[14] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_invx05 \SADR/MAINSADR/U349  ( .ZN(\SADR/MAINSADR/n8807 ), .A(
        \SADR/operand[10] ) );
    snl_muxi21x1 \SADR/MAINSADR/U145  ( .ZN(\pgregadrh[5] ), .A(
        \SADR/MAINSADR/n8769 ), .B(\SADR/MAINSADR/n8748 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U162  ( .ZN(\pgregadrh[18] ), .A(
        \SADR/MAINSADR/n8788 ), .B(\SADR/MAINSADR/n8776 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U252  ( .ZN(\SADR/MAINSADR/n8744 ), .A(
        \SADR/MAINSADR/n8704 ), .B(\SADR/pgaddwxyz[20] ), .C(
        \SADR/MAINSADR/n8706 ), .D(\SADR/pgaddxyz[20] ), .E(
        \SADR/MAINSADR/n8708 ), .F(\SADR/pgaddwyz[20] ), .G(
        \SADR/MAINSADR/n8710 ), .H(\SADR/pgaddwxz[20] ) );
    snl_muxi21x1 \SADR/MAINSADR/U179  ( .ZN(\SADR/MAINSADR/offset[6] ), .A(
        \SADR/MAINSADR/n8807 ), .B(\SADR/MAINSADR/n8808 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi222x0 \SADR/MAINSADR/U275  ( .ZN(\SADR/MAINSADR/n8825 ), .A(
        \pk_indw_h[7] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[7] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[7] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U249  ( .ZN(\SADR/MAINSADR/n8738 ), .A(
        \SADR/pgaddwxy[21] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[21] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[21] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[21] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi012x1 \SADR/MAINSADR/U50  ( .ZN(\SADR/MAINSADR/n8640 ), .A(
        \SADR/MAINSADR/addindoff[20] ), .B(\SADR/MAINSADR/n8638 ), .C(
        \SADR/MAINSADR/n8639 ) );
    snl_muxi21x1 \SADR/MAINSADR/U77  ( .ZN(\SADR/MAINSADR/n8685 ), .A(
        \SADR/MAINSADR/addindoff[3] ), .B(\SADR/m_fadrl[7] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_invx05 \SADR/MAINSADR/U92  ( .ZN(\SADR/MAINSADR/n8649 ), .A(
        \SADR/operand[1] ) );
    snl_nand02x1 \SADR/MAINSADR/U375  ( .ZN(\SADR/MAINSADR/n8755 ), .A(
        \SADR/MAINSADR/oddadd_p1[4] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_and02x1 \SADR/MAINSADR/U117  ( .Z(\SADR/MAINSADR/n8717 ), .A(
        \SADR/MAINSADR/n8709 ), .B(\SADR/MAINSADR/n8707 ) );
    snl_invx05 \SADR/MAINSADR/U352  ( .ZN(\SADR/MAINSADR/n8813 ), .A(
        \SADR/operand[14] ) );
    snl_muxi21x1 \SADR/MAINSADR/U227  ( .ZN(\SADR/MAINSADR/index[16] ), .A(
        \SADR/MAINSADR/n8882 ), .B(\SADR/MAINSADR/n8887 ), .S(ph_lwdsrc_h) );
    snl_muxi21x1 \SADR/MAINSADR/U436  ( .ZN(\pgsdprlh[13] ), .A(
        \SADR/MAINSADR/n8683 ), .B(\SADR/MAINSADR/n8693 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_muxi21x1 \SADR/MAINSADR/U200  ( .ZN(\SADR/MAINSADR/index[8] ), .A(
        \SADR/MAINSADR/n8819 ), .B(\SADR/MAINSADR/n8824 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U390  ( .ZN(\SADR/MAINSADR/n8801 ), .A(
        \SADR/MAINSADR/oddadd_p1[10] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_muxi21x1 \SADR/MAINSADR/U411  ( .ZN(\pgsdprlh[9] ), .A(
        \SADR/MAINSADR/n8682 ), .B(\SADR/MAINSADR/n8683 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_oai012x1 \SADR/MAINSADR/U58  ( .ZN(\pgsdprlh[0] ), .A(
        \SADR/MAINSADR/n8635 ), .B(\SADR/MAINSADR/n8647 ), .C(
        \SADR/MAINSADR/n8648 ) );
    snl_invx05 \SADR/MAINSADR/U130  ( .ZN(\SADR/MAINSADR/n8645 ), .A(
        \SADR/operand[21] ) );
    snl_oa112x1 \SADR/MAINSADR/U138  ( .Z(\SADR/MAINSADR/n8757 ), .A(
        \SADR/MAINSADR/n8678 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8758 ), .D(\SADR/MAINSADR/n8759 ) );
    snl_muxi21x1 \SADR/MAINSADR/U194  ( .ZN(\SADR/MAINSADR/offset[10] ), .A(
        \SADR/MAINSADR/n8813 ), .B(\SADR/MAINSADR/n8807 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi222x0 \SADR/MAINSADR/U283  ( .ZN(\SADR/MAINSADR/n8835 ), .A(
        \pk_indw_h[5] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[5] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[5] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U313  ( .ZN(\SADR/MAINSADR/n8880 ), .A(
        \SADR/pgaddwxy[17] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[17] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[17] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[17] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U334  ( .ZN(\SADR/MAINSADR/n8904 ), .A(
        \SADR/pgaddwz[12] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[12] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[12] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[12] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U208  ( .ZN(\SADR/MAINSADR/index[4] ), .A(
        \SADR/MAINSADR/n8839 ), .B(\SADR/MAINSADR/n8844 ), .S(ph_lwdsrc_h) );
    snl_nand23x1 \SADR/MAINSADR/U398  ( .ZN(\SADR/MAINSADR/n8922 ), .A(
        \SADR/MAINSADR/n8921 ), .B(\SADR/MAINSADR/n8920 ), .C(ph_wrdsrc_h) );
    snl_muxi21x1 \SADR/MAINSADR/U419  ( .ZN(\pgsdprlh[5] ), .A(
        \SADR/MAINSADR/n8687 ), .B(\SADR/MAINSADR/n8682 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi222x0 \SADR/MAINSADR/U16  ( .ZN(\SADR/MAINSADR/n8672 ), .A(
        \SADR/MAINSADR/oddadd_m1[21] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[20] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[20] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U18  ( .ZN(\SADR/MAINSADR/n8775 ), .A(
        \SADR/MAINSADR/oddadd_m1[19] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[18] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[18] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_invx1 \SADR/MAINSADR/U36  ( .ZN(\SADR/MAINSADR/n8918 ), .A(
        \SADR/MAINSADR/n8661 ) );
    snl_oa112x1 \SADR/MAINSADR/U156  ( .Z(\SADR/MAINSADR/n8782 ), .A(
        \SADR/MAINSADR/n8690 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8783 ), .D(\SADR/MAINSADR/n8784 ) );
    snl_muxi21x1 \SADR/MAINSADR/U171  ( .ZN(\pgregadrh[13] ), .A(
        \SADR/MAINSADR/n8745 ), .B(\SADR/MAINSADR/n8791 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U241  ( .ZN(\SADR/MAINSADR/n8728 ), .A(
        \SADR/pgaddwxy[23] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[23] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[23] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[23] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U266  ( .ZN(\SADR/MAINSADR/n8816 ), .A(
        \SADR/pgaddwz[9] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[9] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[9] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[9] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_nor02x2 \SADR/MAINSADR/U43  ( .ZN(\SADR/MAINSADR/n8676 ), .A(
        \SADR/MAINSADR/n8694 ), .B(\SADR/MAINSADR/n8655 ) );
    snl_aoib122x0 \SADR/MAINSADR/U64  ( .ZN(\SADR/MAINSADR/n8665 ), .A(
        \SADR/MAINSADR/n8666 ), .B(\SADR/MAINSADR/oddadd[23] ), .C(
        \SADR/MAINSADR/oddadd_p1[23] ), .D(\SADR/MAINSADR/n8667 ), .E(
        \SADR/MAINSADR/n8668 ) );
    snl_muxi21x1 \SADR/MAINSADR/U81  ( .ZN(\SADR/MAINSADR/n8688 ), .A(
        \SADR/MAINSADR/addindoff[18] ), .B(\SADR/m_fadrl[22] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U341  ( .ZN(\SADR/MAINSADR/n8915 ), .A(
        \SADR/pgaddwxy[10] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[10] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[10] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[10] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_and02x1 \SADR/MAINSADR/U366  ( .Z(\SADR/MAINSADR/n8639 ), .A(
        \SADR/m_fadrl[23] ), .B(\SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U104  ( .Z(\SADR/MAINSADR/n8704 ), .A(
        \SADR/MAINSADR/n8703 ), .B(\SADR/MAINSADR/n8702 ) );
    snl_and04x1 \SADR/MAINSADR/U234  ( .Z(\SADR/MAINSADR/n8907 ), .A(
        \SADR/MAINSADR/n8908 ), .B(\SADR/MAINSADR/n8909 ), .C(
        \SADR/MAINSADR/n8910 ), .D(\SADR/MAINSADR/n8911 ) );
    snl_invx05 \SADR/MAINSADR/U425  ( .ZN(\SADR/MAINSADR/oddadd[17] ), .A(
        \SADR/MAINSADR/n8689 ) );
    snl_aoi012x1 \SADR/MAINSADR/U51  ( .ZN(\SADR/MAINSADR/n8641 ), .A(
        \SADR/MAINSADR/addindoff[21] ), .B(\SADR/MAINSADR/n8638 ), .C(
        \SADR/MAINSADR/n8639 ) );
    snl_muxi21x1 \SADR/MAINSADR/U76  ( .ZN(\SADR/MAINSADR/n8684 ), .A(
        \SADR/MAINSADR/addindoff[4] ), .B(\SADR/m_fadrl[8] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U116  ( .Z(\SADR/MAINSADR/n8716 ), .A(
        \SADR/MAINSADR/n8711 ), .B(\SADR/MAINSADR/n8705 ) );
    snl_and02x1 \SADR/MAINSADR/U123  ( .Z(\SADR/MAINSADR/n8723 ), .A(
        \SADR/MAINSADR/n8719 ), .B(\SADR/MAINSADR/n8705 ) );
    snl_muxi21x1 \SADR/MAINSADR/U213  ( .ZN(\SADR/MAINSADR/index[23] ), .A(
        \SADR/MAINSADR/n8859 ), .B(\SADR/MAINSADR/n8860 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U383  ( .ZN(\SADR/MAINSADR/n8780 ), .A(
        \SADR/MAINSADR/oddadd_p1[17] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_muxi21x1 \SADR/MAINSADR/U402  ( .ZN(\pgsdprlh[12] ), .A(
        \SADR/MAINSADR/n8675 ), .B(\SADR/MAINSADR/n8677 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U298  ( .ZN(\SADR/MAINSADR/n8856 ), .A(
        \SADR/pgaddwz[1] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[1] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[1] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[1] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U308  ( .ZN(\SADR/MAINSADR/n8876 ), .A(
        \SADR/pgaddwxyz[18] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[18] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[18] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[18] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_and04x1 \SADR/MAINSADR/U226  ( .Z(\SADR/MAINSADR/n8887 ), .A(
        \SADR/MAINSADR/n8888 ), .B(\SADR/MAINSADR/n8889 ), .C(
        \SADR/MAINSADR/n8890 ), .D(\SADR/MAINSADR/n8891 ) );
    snl_invx05 \SADR/MAINSADR/U131  ( .ZN(\SADR/MAINSADR/n8644 ), .A(
        \SADR/operand[20] ) );
    snl_and04x1 \SADR/MAINSADR/U201  ( .Z(\SADR/MAINSADR/n8829 ), .A(
        \SADR/MAINSADR/n8830 ), .B(\SADR/MAINSADR/n8831 ), .C(
        \SADR/MAINSADR/n8832 ), .D(\SADR/MAINSADR/n8833 ) );
    snl_invx05 \SADR/MAINSADR/U391  ( .ZN(\SADR/MAINSADR/n8862 ), .A(
        \SADR/MAINSADR/n8740 ) );
    snl_invx05 \SADR/MAINSADR/U410  ( .ZN(\SADR/MAINSADR/oddadd[5] ), .A(
        \SADR/MAINSADR/n8682 ) );
    snl_mux21x1 \SADR/MAINSADR/U178  ( .Z(\SADR/MAINSADR/offset[7] ), .A(
        \SADR/operand[11] ), .B(\SADR/operand[7] ), .S(\SADR/MAINSADR/n8635 )
         );
    snl_aoi222x0 \SADR/MAINSADR/U23  ( .ZN(\SADR/MAINSADR/n8790 ), .A(
        \SADR/MAINSADR/oddadd_m1[14] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[13] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[13] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_aoi222x0 \SADR/MAINSADR/U24  ( .ZN(\SADR/MAINSADR/n8793 ), .A(
        \SADR/MAINSADR/oddadd_m1[13] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[12] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[12] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_invx05 \SADR/MAINSADR/U88  ( .ZN(\SADR/MAINSADR/n8694 ), .A(
        ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U93  ( .ZN(\SADR/MAINSADR/n8647 ), .A(
        \SADR/operand[0] ) );
    snl_aoi2222x0 \SADR/MAINSADR/U248  ( .ZN(\SADR/MAINSADR/n8739 ), .A(
        \SADR/pgaddwxyz[21] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[21] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[21] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[21] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_invx05 \SADR/MAINSADR/U353  ( .ZN(\SADR/MAINSADR/n8812 ), .A(
        \SADR/operand[16] ) );
    snl_nand02x1 \SADR/MAINSADR/U374  ( .ZN(\SADR/MAINSADR/n8746 ), .A(
        \SADR/MAINSADR/oddadd_p1[9] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_oa112x1 \SADR/MAINSADR/U144  ( .Z(\SADR/MAINSADR/n8769 ), .A(
        \SADR/MAINSADR/n8687 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8770 ), .D(\SADR/MAINSADR/n8771 ) );
    snl_oa112x1 \SADR/MAINSADR/U163  ( .Z(\SADR/MAINSADR/n8791 ), .A(
        \SADR/MAINSADR/n8693 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8792 ), .D(\SADR/MAINSADR/n8793 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U253  ( .ZN(\SADR/MAINSADR/n8743 ), .A(
        \SADR/MAINSADR/n8712 ), .B(\SADR/pgaddwxy[20] ), .C(
        \SADR/MAINSADR/n8714 ), .D(\SADR/pgaddyz[20] ), .E(
        \SADR/MAINSADR/n8715 ), .F(\SADR/pgaddxz[20] ), .G(
        \SADR/MAINSADR/n8716 ), .H(\SADR/pgaddxy[20] ) );
    snl_invx05 \SADR/MAINSADR/U348  ( .ZN(\SADR/MAINSADR/n8804 ), .A(
        \SADR/operand[9] ) );
    snl_aoi2222x0 \SADR/MAINSADR/U274  ( .ZN(\SADR/MAINSADR/n8826 ), .A(
        \SADR/pgaddwz[7] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[7] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[7] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[7] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U181  ( .ZN(\SADR/MAINSADR/offset[4] ), .A(
        \SADR/MAINSADR/n8806 ), .B(\SADR/MAINSADR/n8695 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_muxi21x1 \SADR/MAINSADR/U186  ( .ZN(\SADR/MAINSADR/offset[18] ), .A(
        \SADR/MAINSADR/n8646 ), .B(\SADR/MAINSADR/n8810 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi222x0 \SADR/MAINSADR/U291  ( .ZN(\SADR/MAINSADR/n8845 ), .A(
        \pk_indw_h[3] ), .B(\SADR/MAINSADR/n8724 ), .C(\pk_indy_h[3] ), .D(
        \SADR/MAINSADR/n8722 ), .E(\pk_indx_h[3] ), .F(\SADR/MAINSADR/n8723 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U301  ( .ZN(\SADR/MAINSADR/n8866 ), .A(
        \SADR/pgaddwxy[19] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[19] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[19] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[19] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U326  ( .ZN(\SADR/MAINSADR/n8894 ), .A(
        \SADR/pgaddwz[14] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[14] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[14] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[14] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U296  ( .ZN(\SADR/MAINSADR/n8858 ), .A(
        \SADR/pgaddwxyz[1] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[1] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[1] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[1] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U306  ( .ZN(\SADR/MAINSADR/n8869 ), .A(
        \SADR/pgaddwz[0] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[0] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[0] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[0] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U321  ( .ZN(\SADR/MAINSADR/n8890 ), .A(
        \SADR/pgaddwxy[15] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[15] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[15] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[15] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_invx05 \SADR/MAINSADR/U368  ( .ZN(\SADR/MAINSADR/oddadd[19] ), .A(
        \SADR/MAINSADR/n8637 ) );
    snl_aoi222x0 \SADR/MAINSADR/U31  ( .ZN(\SADR/MAINSADR/n8762 ), .A(
        \SADR/MAINSADR/oddadd_m1[3] ), .B(\SADR/MAINSADR/n8698 ), .C(
        \SADR/MAINSADR/oddadd_m2[2] ), .D(\SADR/MAINSADR/n8917 ), .E(
        \SADR/MAINSADR/oddadd_p2[2] ), .F(\SADR/MAINSADR/n8918 ) );
    snl_invx2 \SADR/MAINSADR/U38  ( .ZN(\SADR/MAINSADR/n8634 ), .A(
        \SADR/MAINSADR/n8633 ) );
    snl_muxi21x1 \SADR/MAINSADR/U143  ( .ZN(\pgregadrh[6] ), .A(
        \SADR/MAINSADR/n8766 ), .B(\SADR/MAINSADR/n8763 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U273  ( .ZN(\SADR/MAINSADR/n8827 ), .A(
        \SADR/pgaddwxy[7] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[7] ), 
        .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[7] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[7] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_muxi21x1 \SADR/MAINSADR/U158  ( .ZN(\pgregadrh[1] ), .A(
        \SADR/MAINSADR/n8649 ), .B(\SADR/MAINSADR/n8769 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_muxi21x1 \SADR/MAINSADR/U164  ( .ZN(\pgregadrh[17] ), .A(
        \SADR/MAINSADR/n8791 ), .B(\SADR/MAINSADR/n8779 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U254  ( .ZN(\SADR/MAINSADR/n8742 ), .A(
        \SADR/MAINSADR/n8717 ), .B(\SADR/pgaddwz[20] ), .C(
        \SADR/MAINSADR/n8718 ), .D(\SADR/pgaddwy[20] ), .E(
        \SADR/MAINSADR/n8720 ), .F(\SADR/pgaddwx[20] ), .G(
        \SADR/MAINSADR/n8721 ), .H(\pk_indz_h[20] ) );
    snl_aoi2222x0 \SADR/MAINSADR/U268  ( .ZN(\SADR/MAINSADR/n8823 ), .A(
        \SADR/pgaddwxyz[8] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[8] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[8] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[8] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_oai012x2 \SADR/MAINSADR/U44  ( .ZN(\SADR/MAINSADR/n8667 ), .A(
        ph_lwdsrc_h), .B(\SADR/MAINSADR/n8697 ), .C(\SADR/MAINSADR/n8699 ) );
    snl_nor02x1 \SADR/MAINSADR/U56  ( .ZN(\SADR/MAINSADR/offset[22] ), .A(
        \SADR/MAINSADR/n8643 ), .B(\SADR/MAINSADR/n8646 ) );
    snl_invx05 \SADR/MAINSADR/U94  ( .ZN(\SADR/MAINSADR/n8695 ), .A(
        \SADR/operand[4] ) );
    snl_oa112x1 \SADR/MAINSADR/U136  ( .Z(\SADR/MAINSADR/n8754 ), .A(
        \SADR/MAINSADR/n8684 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8755 ), .D(\SADR/MAINSADR/n8756 ) );
    snl_invx05 \SADR/MAINSADR/U354  ( .ZN(\SADR/MAINSADR/n8811 ), .A(
        \SADR/operand[17] ) );
    snl_nand02x1 \SADR/MAINSADR/U373  ( .ZN(\SADR/MAINSADR/n8749 ), .A(
        \SADR/MAINSADR/oddadd_p1[5] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_muxi21x1 \SADR/MAINSADR/U206  ( .ZN(\SADR/MAINSADR/index[5] ), .A(
        \SADR/MAINSADR/n8834 ), .B(\SADR/MAINSADR/n8839 ), .S(ph_lwdsrc_h) );
    snl_nand04x0 \SADR/MAINSADR/U396  ( .ZN(\SADR/MAINSADR/n8923 ), .A(
        \SADR/MAINSADR/n8642 ), .B(\SADR/MAINSADR/n8641 ), .C(
        \SADR/MAINSADR/n8640 ), .D(\SADR/MAINSADR/n8637 ) );
    snl_muxi21x1 \SADR/MAINSADR/U417  ( .ZN(\pgsdprlh[6] ), .A(
        \SADR/MAINSADR/n8686 ), .B(\SADR/MAINSADR/n8680 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U71  ( .ZN(\SADR/MAINSADR/n8679 ), .A(
        \SADR/MAINSADR/addindoff[11] ), .B(\SADR/m_fadrl[15] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_muxi21x1 \SADR/MAINSADR/U221  ( .ZN(\SADR/MAINSADR/index[19] ), .A(
        \SADR/MAINSADR/n8863 ), .B(\SADR/MAINSADR/n8872 ), .S(ph_lwdsrc_h) );
    snl_invx05 \SADR/MAINSADR/U430  ( .ZN(\SADR/MAINSADR/oddadd[14] ), .A(
        \SADR/MAINSADR/n8692 ) );
    snl_nor02x1 \SADR/MAINSADR/U111  ( .ZN(\SADR/MAINSADR/n8711 ), .A(
        \SADR/MAINSADR/n8701 ), .B(\SADR/operand[24] ) );
    snl_and02x1 \SADR/MAINSADR/U124  ( .Z(\SADR/MAINSADR/n8724 ), .A(
        \SADR/MAINSADR/n8719 ), .B(\SADR/MAINSADR/n8707 ) );
    snl_muxi21x1 \SADR/MAINSADR/U214  ( .ZN(\SADR/MAINSADR/index[22] ), .A(
        \SADR/MAINSADR/n8860 ), .B(\SADR/MAINSADR/n8861 ), .S(ph_lwdsrc_h) );
    snl_nand02x1 \SADR/MAINSADR/U384  ( .ZN(\SADR/MAINSADR/n8783 ), .A(
        \SADR/MAINSADR/oddadd_p1[16] ), .B(\SADR/MAINSADR/n8667 ) );
    snl_muxi21x1 \SADR/MAINSADR/U405  ( .ZN(\pgsdprlh[11] ), .A(
        \SADR/MAINSADR/n8678 ), .B(\SADR/MAINSADR/n8679 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi013x0 \SADR/MAINSADR/U63  ( .ZN(\SADR/MAINSADR/n8660 ), .A(
        \SADR/MAINSADR/n8661 ), .B(\SADR/MAINSADR/n8662 ), .C(
        \SADR/MAINSADR/n8663 ), .D(\SADR/MAINSADR/n8664 ) );
    snl_muxi21x1 \SADR/MAINSADR/U233  ( .ZN(\SADR/MAINSADR/index[13] ), .A(
        \SADR/MAINSADR/n8897 ), .B(\SADR/MAINSADR/n8902 ), .S(ph_lwdsrc_h) );
    snl_mux21x1 \SADR/MAINSADR/U422  ( .Z(\pgsdprlh[23] ), .A(
        \SADR/MAINSADR/oddadd[19] ), .B(\SADR/MAINSADR/oddadd[23] ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_muxi21x1 \SADR/MAINSADR/U86  ( .ZN(\SADR/MAINSADR/n8693 ), .A(
        \SADR/MAINSADR/addindoff[13] ), .B(\SADR/m_fadrl[17] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U103  ( .Z(\SADR/MAINSADR/n8703 ), .A(
        \SADR/operand[27] ), .B(\SADR/operand[26] ) );
    snl_muxi21x1 \SADR/MAINSADR/U188  ( .ZN(\SADR/MAINSADR/offset[16] ), .A(
        \SADR/MAINSADR/n8644 ), .B(\SADR/MAINSADR/n8812 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U328  ( .ZN(\SADR/MAINSADR/n8901 ), .A(
        \SADR/pgaddwxyz[13] ), .B(\SADR/MAINSADR/n8704 ), .C(
        \SADR/pgaddxyz[13] ), .D(\SADR/MAINSADR/n8706 ), .E(
        \SADR/pgaddwyz[13] ), .F(\SADR/MAINSADR/n8708 ), .G(
        \SADR/pgaddwxz[13] ), .H(\SADR/MAINSADR/n8710 ) );
    snl_invx05 \SADR/MAINSADR/U346  ( .ZN(\SADR/MAINSADR/n8808 ), .A(
        \SADR/operand[6] ) );
    snl_invx05 \SADR/MAINSADR/U361  ( .ZN(\SADR/intbitno[2] ), .A(
        \SADR/MAINSADR/n8652 ) );
    snl_muxi21x1 \SADR/MAINSADR/U151  ( .ZN(\pgregadrh[23] ), .A(
        \SADR/MAINSADR/n8773 ), .B(\SADR/MAINSADR/n8665 ), .S(
        \SADR/MAINSADR/n8635 ) );
    snl_aoi022x1 \SADR/MAINSADR/U261  ( .ZN(\SADR/MAINSADR/n8926 ), .A(
        \SADR/pgovfxz ), .B(\SADR/MAINSADR/n8715 ), .C(\SADR/pgovfxy ), .D(
        \SADR/MAINSADR/n8716 ) );
    snl_muxi21x1 \SADR/MAINSADR/U176  ( .ZN(\SADR/MAINSADR/offset[9] ), .A(
        \SADR/MAINSADR/n8803 ), .B(\SADR/MAINSADR/n8804 ), .S(
        \SADR/MAINSADR/n8634 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U246  ( .ZN(\SADR/MAINSADR/n8732 ), .A(
        \SADR/pgaddwz[22] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[22] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[22] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[22] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_muxi21x1 \SADR/MAINSADR/U78  ( .ZN(\SADR/MAINSADR/n8686 ), .A(
        \SADR/MAINSADR/addindoff[2] ), .B(\SADR/m_fadrl[6] ), .S(
        \SADR/MAINSADR/n8676 ) );
    snl_and02x1 \SADR/MAINSADR/U118  ( .Z(\SADR/MAINSADR/n8718 ), .A(
        \SADR/MAINSADR/n8711 ), .B(\SADR/MAINSADR/n8707 ) );
    snl_mux21x1 \SADR/MAINSADR/U193  ( .Z(\SADR/MAINSADR/offset[11] ), .A(
        \SADR/operand[15] ), .B(\SADR/operand[11] ), .S(\SADR/MAINSADR/n8635 )
         );
    snl_aoi2222x0 \SADR/MAINSADR/U284  ( .ZN(\SADR/MAINSADR/n8843 ), .A(
        \SADR/pgaddwxyz[4] ), .B(\SADR/MAINSADR/n8704 ), .C(\SADR/pgaddxyz[4] 
        ), .D(\SADR/MAINSADR/n8706 ), .E(\SADR/pgaddwyz[4] ), .F(
        \SADR/MAINSADR/n8708 ), .G(\SADR/pgaddwxz[4] ), .H(
        \SADR/MAINSADR/n8710 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U333  ( .ZN(\SADR/MAINSADR/n8905 ), .A(
        \SADR/pgaddwxy[12] ), .B(\SADR/MAINSADR/n8712 ), .C(\SADR/pgaddyz[12] 
        ), .D(\SADR/MAINSADR/n8714 ), .E(\SADR/pgaddxz[12] ), .F(
        \SADR/MAINSADR/n8715 ), .G(\SADR/pgaddxy[12] ), .H(
        \SADR/MAINSADR/n8716 ) );
    snl_aoi2222x0 \SADR/MAINSADR/U314  ( .ZN(\SADR/MAINSADR/n8879 ), .A(
        \SADR/pgaddwz[17] ), .B(\SADR/MAINSADR/n8717 ), .C(\SADR/pgaddwy[17] ), 
        .D(\SADR/MAINSADR/n8718 ), .E(\SADR/pgaddwx[17] ), .F(
        \SADR/MAINSADR/n8720 ), .G(\pk_indz_h[17] ), .H(\SADR/MAINSADR/n8721 )
         );
    snl_and04x1 \SADR/MAINSADR/U228  ( .Z(\SADR/MAINSADR/n8892 ), .A(
        \SADR/MAINSADR/n8893 ), .B(\SADR/MAINSADR/n8894 ), .C(
        \SADR/MAINSADR/n8895 ), .D(\SADR/MAINSADR/n8896 ) );
    snl_ao022x1 \REGF/pbmemff21/U134  ( .Z(\REGF/pbmemff21/RO_PC19B72[12] ), 
        .A(PDLIN[12]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[12] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U141  ( .Z(\REGF/pbmemff21/RO_PPC19B114[2] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[2] ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[15]  ( .Q(\pk_pc_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[15] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_bufx2 \REGF/pbmemff21/U115  ( .Z(\REGF/pbmemff21/n6969 ), .A(
        \REGF/n8052 ) );
    snl_ao022x4 \REGF/pbmemff21/U120  ( .Z(\REGF/pbmemff21/RO_PC19B72[17] ), 
        .A(PDLIN[17]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[17] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_ao022x4 \REGF/pbmemff21/U121  ( .Z(\REGF/pbmemff21/RO_PC19B72[7] ), 
        .A(PDLIN[7]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[7] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_ao022x1 \REGF/pbmemff21/U126  ( .Z(\REGF/pbmemff21/RO_PC19B72[1] ), 
        .A(PDLIN[1]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[1] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U148  ( .Z(\REGF/pbmemff21/RO_PPC19B114[9] ), 
        .A(\pk_pc_h[9] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_and02x1 \REGF/pbmemff21/U153  ( .Z(\REGF/pbmemff21/RO_PPC19B114[14] ), 
        .A(\pk_pc_h[14] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[11]  ( .Q(\pk_pc_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[11] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[18]  ( .Q(\pk_pc_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[18] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U128  ( .Z(\REGF/pbmemff21/RO_PC19B72[3] ), 
        .A(PDLIN[3]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[3] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U154  ( .Z(\REGF/pbmemff21/RO_PPC19B114[15] ), 
        .A(\pk_pc_h[15] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[13]  ( .Q(\pk_pc_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[13] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U133  ( .Z(\REGF/pbmemff21/RO_PC19B72[11] ), 
        .A(PDLIN[11]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[11] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U146  ( .Z(\REGF/pbmemff21/RO_PPC19B114[7] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[7] ) );
    snl_and02x1 \REGF/pbmemff21/U155  ( .Z(\REGF/pbmemff21/RO_PPC19B114[16] ), 
        .A(\pk_pc_h[16] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[17]  ( .Q(\pk_pc_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[17] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[4]  ( .Q(\REGF/RO_PPCN[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[4] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[5]  ( .Q(\pk_pc_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[5] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[13]  ( .Q(\REGF/RO_PPCN[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[13] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U132  ( .Z(\REGF/pbmemff21/RO_PC19B72[10] ), 
        .A(PDLIN[10]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[10] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_nand12x2 \REGF/pbmemff21/U116  ( .ZN(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .A(polcore_end), .B(
        \REGF/pbmemff21/n6970 ) );
    snl_nor02x4 \REGF/pbmemff21/U117  ( .ZN(\REGF/pbmemff21/n6970 ), .A(
        \pk_rwrit_h[44] ), .B(\pk_rwrit_h[59] ) );
    snl_ao022x4 \REGF/pbmemff21/U119  ( .Z(\REGF/pbmemff21/RO_PC19B72[8] ), 
        .A(PDLIN[8]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[8] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_ao022x1 \REGF/pbmemff21/U127  ( .Z(\REGF/pbmemff21/RO_PC19B72[2] ), 
        .A(PDLIN[2]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[2] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_ao022x1 \REGF/pbmemff21/U129  ( .Z(\REGF/pbmemff21/RO_PC19B72[4] ), 
        .A(PDLIN[4]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[4] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U147  ( .Z(\REGF/pbmemff21/RO_PPC19B114[8] ), 
        .A(\pk_pc_h[8] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[8]  ( .Q(\pk_pc_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[8] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[0]  ( .Q(\REGF/RO_PPCN[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[0] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[1]  ( .Q(\pk_pc_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[1] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[17]  ( .Q(\REGF/RO_PPCN[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[17] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[9]  ( .Q(\REGF/RO_PPCN[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[9] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U135  ( .Z(\REGF/pbmemff21/RO_PC19B72[13] ), 
        .A(PDLIN[13]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[13] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U140  ( .Z(\REGF/pbmemff21/RO_PPC19B114[1] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[1] ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[3]  ( .Q(\pk_pc_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[3] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[15]  ( .Q(\REGF/RO_PPCN[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[15] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[2]  ( .Q(\REGF/RO_PPCN[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[2] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[11]  ( .Q(\REGF/RO_PPCN[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[11] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U137  ( .Z(\REGF/pbmemff21/RO_PC19B72[16] ), 
        .A(PDLIN[16]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[16] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U149  ( .Z(\REGF/pbmemff21/RO_PPC19B114[10] ), 
        .A(\pk_pc_h[10] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_and02x1 \REGF/pbmemff21/U152  ( .Z(\REGF/pbmemff21/RO_PPC19B114[13] ), 
        .A(\pk_pc_h[13] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[7]  ( .Q(\pk_pc_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[7] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[6]  ( .Q(\REGF/RO_PPCN[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[6] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[18]  ( .Q(\REGF/RO_PPCN[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[18] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff21/U142  ( .Z(\REGF/pbmemff21/RO_PPC19B114[3] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[3] ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[6]  ( .Q(\pk_pc_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[6] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[10]  ( .Q(\REGF/RO_PPCN[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[10] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[7]  ( .Q(\REGF/RO_PPCN[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[7] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_ao022x4 \REGF/pbmemff21/U122  ( .Z(\REGF/pbmemff21/RO_PC19B72[15] ), 
        .A(PDLIN[15]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[15] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_ao022x1 \REGF/pbmemff21/U125  ( .Z(\REGF/pbmemff21/RO_PC19B72[0] ), 
        .A(PDLIN[0]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[0] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U150  ( .Z(\REGF/pbmemff21/RO_PPC19B114[11] ), 
        .A(\pk_pc_h[11] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[2]  ( .Q(\pk_pc_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[2] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[14]  ( .Q(\REGF/RO_PPCN[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[14] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[3]  ( .Q(\REGF/RO_PPCN[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[3] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff21/U139  ( .Z(\REGF/pbmemff21/RO_PPC19B114[0] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[0] ) );
    snl_and02x1 \REGF/pbmemff21/U157  ( .Z(\REGF/pbmemff21/RO_PPC19B114[18] ), 
        .A(\pk_pc_h[18] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[9]  ( .Q(\pk_pc_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[9] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[16]  ( .Q(\REGF/RO_PPCN[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[16] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[1]  ( .Q(\REGF/RO_PPCN[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[1] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[8]  ( .Q(\REGF/RO_PPCN[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[8] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff21/U145  ( .Z(\REGF/pbmemff21/RO_PPC19B114[6] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[6] ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[0]  ( .Q(\pk_pc_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[0] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[5]  ( .Q(\REGF/RO_PPCN[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[5] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[4]  ( .Q(\pk_pc_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[4] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_and08x1 \REGF/pbmemff21/U123  ( .Z(pk_pcovf_h), .A(\pk_pc_h[0] ), .B(
        \pk_pc_h[1] ), .C(\pk_pc_h[2] ), .D(\pk_pc_h[3] ), .E(\pk_pc_h[4] ), 
        .F(\pk_pc_h[5] ), .G(\pk_pc_h[6] ), .H(\pk_pc_h[7] ) );
    snl_ao022x1 \REGF/pbmemff21/U130  ( .Z(\REGF/pbmemff21/RO_PC19B72[5] ), 
        .A(PDLIN[5]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[5] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PPC19B_reg[12]  ( .Q(\REGF/RO_PPCN[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PPC19B114[12] ), .SE(\REGF/pbmemff21/n_853 ), .CP(
        SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U138  ( .Z(\REGF/pbmemff21/RO_PC19B72[18] ), 
        .A(PDLIN[18]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[18] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U156  ( .Z(\REGF/pbmemff21/RO_PPC19B114[17] ), 
        .A(\pk_pc_h[17] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[16]  ( .Q(\pk_pc_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[16] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_ao022x1 \REGF/pbmemff21/U131  ( .Z(\REGF/pbmemff21/RO_PC19B72[6] ), 
        .A(PDLIN[6]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[6] ), 
        .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U144  ( .Z(\REGF/pbmemff21/RO_PPC19B114[5] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[5] ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[12]  ( .Q(\pk_pc_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[12] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_ao022x4 \REGF/pbmemff21/U118  ( .Z(\REGF/pbmemff21/RO_PC19B72[9] ), 
        .A(\pk_rwrit_h[59] ), .B(PDLIN[9]), .C(\REGF/pbmemff21/n6970 ), .D(
        \REGF/pbmemff21/RO_PC19BT[9] ) );
    snl_ao012x1 \REGF/pbmemff21/U124  ( .Z(\REGF/pbmemff21/n_853 ), .A(
        polcore_end), .B(\pk_rread_h[50] ), .C(\pk_rwrit_h[44] ) );
    snl_ao022x1 \REGF/pbmemff21/U136  ( .Z(\REGF/pbmemff21/RO_PC19B72[14] ), 
        .A(PDLIN[14]), .B(\pk_rwrit_h[59] ), .C(\REGF/pbmemff21/RO_PC19BT[14] 
        ), .D(\REGF/pbmemff21/n6970 ) );
    snl_and02x1 \REGF/pbmemff21/U143  ( .Z(\REGF/pbmemff21/RO_PPC19B114[4] ), 
        .A(\REGF/pbmemff21/n6971 ), .B(\pk_pc_h[4] ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[10]  ( .Q(\pk_pc_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[10] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \REGF/pbmemff21/U158  ( .ZN(\REGF/pbmemff21/n6971 ), .A(
        \pk_rwrit_h[44] ) );
    snl_and02x1 \REGF/pbmemff21/U151  ( .Z(\REGF/pbmemff21/RO_PPC19B114[12] ), 
        .A(\pk_pc_h[12] ), .B(\REGF/pbmemff21/n6971 ) );
    snl_sffqenrnx1 \REGF/pbmemff21/RO_PC19B_reg[14]  ( .Q(\pk_pc_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff21/n6969 ), .SD(
        \REGF/pbmemff21/RO_PC19B72[14] ), .SE(
        \REGF/pbmemff21/*cell*5483/U4/CONTROL1 ), .CP(SCLK) );
    snl_nand12x1 \REG_2/ph8dec_1/U6  ( .ZN(\REG_2/ncnt1[2] ), .A(ph_tirtendh), 
        .B(\REG_2/ph8dec_1/n22 ) );
    snl_invx05 \REG_2/ph8dec_1/U7  ( .ZN(\REG_2/ncnt1[0] ), .A(
        \REG_2/RETCNT[0] ) );
    snl_aoi022x1 \REG_2/ph8dec_1/U8  ( .ZN(\REG_2/ncnt1[1] ), .A(
        \REG_2/RETCNT[1] ), .B(\REG_2/ncnt1[0] ), .C(\REG_2/ph8dec_1/n23 ), 
        .D(\REG_2/RETCNT[0] ) );
    snl_nor03x0 \REG_2/ph8dec_1/U9  ( .ZN(ph_tirtendh), .A(\REG_2/RETCNT[0] ), 
        .B(\REG_2/RETCNT[2] ), .C(\REG_2/RETCNT[1] ) );
    snl_oai012x1 \REG_2/ph8dec_1/U10  ( .ZN(\REG_2/ph8dec_1/n22 ), .A(
        \REG_2/RETCNT[1] ), .B(\REG_2/RETCNT[0] ), .C(\REG_2/RETCNT[2] ) );
    snl_invx05 \REG_2/ph8dec_1/U11  ( .ZN(\REG_2/ph8dec_1/n23 ), .A(
        \REG_2/RETCNT[1] ) );
    snl_or02x1 \SADR/ADDIDX/U7  ( .Z(\SADR/pgovfwxz ), .A(\SADR/pgovfxz ), .B(
        \SADR/ADDIDX/pgovfwxzT ) );
    snl_or02x1 \SADR/ADDIDX/U8  ( .Z(\SADR/pgovfwxy ), .A(\SADR/pgovfwx ), .B(
        \SADR/ADDIDX/pgovfwxyT ) );
    snl_or02x1 \SADR/ADDIDX/U9  ( .Z(\SADR/pgovfxyz ), .A(\SADR/pgovfyz ), .B(
        \SADR/ADDIDX/pgovfxyzT ) );
    snl_or02x1 \SADR/ADDIDX/U10  ( .Z(\SADR/pgovfwyz ), .A(\SADR/pgovfwy ), 
        .B(\SADR/ADDIDX/pgovfwyzT ) );
    snl_or03x1 \SADR/ADDIDX/U11  ( .Z(\SADR/pgovfwxyz ), .A(
        \SADR/ADDIDX/pgovfwxyzT ), .B(\SADR/pgovfwz ), .C(\SADR/pgovfxy ) );
    snl_oai2222x0 \SAEXE/SRC2/U94  ( .ZN(\SAEXE/SRC2/nqst[0] ), .A(
        \SAEXE/seq_end ), .B(\SAEXE/SRC2/n184 ), .C(\SAEXE/singlen ), .D(
        \SAEXE/SRC2/n185 ), .E(pgadrovfh), .F(\SAEXE/SRC2/n186 ), .G(
        \SAEXE/SRC2/eqst[2] ), .H(\SAEXE/SRC2/n187 ) );
    snl_oai112x0 \SAEXE/SRC2/U95  ( .ZN(\SAEXE/SRC2/nqst[1] ), .A(
        \SAEXE/SRC2/n186 ), .B(\SAEXE/SRC2/n188 ), .C(\SAEXE/SRC2/n189 ), .D(
        \SAEXE/SRC2/n190 ) );
    snl_oai112x0 \SAEXE/SRC2/U96  ( .ZN(\SAEXE/SRC2/nqst[2] ), .A(
        \SAEXE/seq_end ), .B(\SAEXE/SRC2/n184 ), .C(\SAEXE/SRC2/n189 ), .D(
        \SAEXE/SRC2/n191 ) );
    snl_and02x1 \SAEXE/SRC2/U113  ( .Z(\SAEXE/SRC2/n206 ), .A(
        \SAEXE/SRC2/eqst[1] ), .B(\SAEXE/SRC2/eqst[2] ) );
    snl_nand03x0 \SAEXE/SRC2/U134  ( .ZN(\SAEXE/SRC2/n220 ), .A(\SAEXE/sequen 
        ), .B(\SAEXE/SRC2/n214 ), .C(\SAEXE/seq_end ) );
    snl_ffqrnx1 \SAEXE/SRC2/eqst_reg[1]  ( .Q(\SAEXE/SRC2/eqst[1] ), .D(
        \SAEXE/SRC2/nqst[1] ), .RN(n10735), .CP(SCLK) );
    snl_oai112x0 \SAEXE/SRC2/U97  ( .ZN(\SAEXE/SRC2/nqst[3] ), .A(
        \SAEXE/SRC2/eqst[2] ), .B(\SAEXE/SRC2/n192 ), .C(\SAEXE/SRC2/n193 ), 
        .D(\SAEXE/SRC2/n194 ) );
    snl_ao2222x1 \SAEXE/SRC2/U98  ( .Z(ph_lblockh), .A(\SAEXE/SRC2/eqst[4] ), 
        .B(\SAEXE/SRC2/n195 ), .C(\SAEXE/SRC2/n196 ), .D(\SAEXE/SRC2/n188 ), 
        .E(\SAEXE/SRC2/n197 ), .F(\SAEXE/SRC2/n198 ), .G(ph_bitsrch), .H(
        \SAEXE/SRC2/n199 ) );
    snl_oai023x0 \SAEXE/SRC2/U101  ( .ZN(\SAEXE/srcwt_st ), .A(
        \SAEXE/SRC2/n203 ), .B(\SAEXE/ph_lber1_h ), .C(\SAEXE/SRC2/n198 ), .D(
        pgadrovfh), .E(\SAEXE/SRC2/n204 ) );
    snl_nor02x1 \SAEXE/SRC2/U108  ( .ZN(\SAEXE/SRC2/n213 ), .A(
        \SAEXE/SRC2/n195 ), .B(\SAEXE/SRC2/eqst[1] ) );
    snl_muxi21x1 \SAEXE/SRC2/U141  ( .ZN(\SAEXE/SRC2/n209 ), .A(
        \SAEXE/SRC2/n215 ), .B(\SAEXE/SRC2/n219 ), .S(\SAEXE/singlen ) );
    snl_nand04x0 \SAEXE/SRC2/U106  ( .ZN(\SAEXE/SRC2/n211 ), .A(
        \SAEXE/srcwrit ), .B(ph_saexe_sth), .C(\SAEXE/singlen ), .D(
        \SAEXE/SRC2/n212 ) );
    snl_and02x1 \SAEXE/SRC2/U121  ( .Z(\SAEXE/SRC2/n218 ), .A(
        \SAEXE/SRC2/n204 ), .B(\SAEXE/SRC2/n216 ) );
    snl_and02x1 \SAEXE/SRC2/U126  ( .Z(\SAEXE/SRC2/n202 ), .A(
        \SAEXE/SRC2/n216 ), .B(\SAEXE/SRC2/n186 ) );
    snl_oai033x0 \SAEXE/SRC2/U99  ( .ZN(\SAEXE/trsc1_h ), .A(\SAEXE/SRC2/n195 
        ), .B(\SAEXE/stage_2nd ), .C(\SAEXE/stage_1st ), .D(\SAEXE/SRC2/n200 ), 
        .E(\SAEXE/SRC2/n201 ), .F(\SAEXE/SRC2/n198 ) );
    snl_nand02x1 \SAEXE/SRC2/U114  ( .ZN(\SAEXE/SRC2/n203 ), .A(
        \SAEXE/SRC2/eqst[4] ), .B(\SAEXE/SRC2/n206 ) );
    snl_nor04x0 \SAEXE/SRC2/U128  ( .ZN(\SAEXE/SRC2/n212 ), .A(
        \SAEXE/SRC2/eqst[2] ), .B(\SAEXE/stage_1st ), .C(\SAEXE/sequen ), .D(
        \SAEXE/srcread ) );
    snl_invx05 \SAEXE/SRC2/U133  ( .ZN(\SAEXE/SRC2/n197 ), .A(
        \SAEXE/SRC2/n203 ) );
    snl_ffqrnx1 \SAEXE/SRC2/eqst_reg[3]  ( .Q(\SAEXE/stage_2nd ), .D(
        \SAEXE/SRC2/nqst[3] ), .RN(n10735), .CP(SCLK) );
    snl_invx05 \SAEXE/SRC2/U107  ( .ZN(\SAEXE/SRC2/n195 ), .A(
        \SAEXE/SRC2/eqst[2] ) );
    snl_oa022x1 \SAEXE/SRC2/U120  ( .Z(\SAEXE/SRC2/n193 ), .A(\SAEXE/seq_end ), 
        .B(\SAEXE/SRC2/n217 ), .C(\SAEXE/SRC2/n207 ), .D(\SAEXE/SRC2/n203 ) );
    snl_nand02x1 \SAEXE/SRC2/U109  ( .ZN(\SAEXE/SRC2/n184 ), .A(
        \SAEXE/SRC2/n213 ), .B(\SAEXE/SRC2/n208 ) );
    snl_nand02x1 \SAEXE/SRC2/U115  ( .ZN(\SAEXE/SRC2/n216 ), .A(
        \SAEXE/SRC2/eqst[4] ), .B(\SAEXE/SRC2/n213 ) );
    snl_invx05 \SAEXE/SRC2/U132  ( .ZN(\SAEXE/SRC2/n196 ), .A(
        \SAEXE/SRC2/n216 ) );
    snl_oa112x1 \SAEXE/SRC2/U129  ( .Z(\SAEXE/SRC2/n194 ), .A(
        \SAEXE/SRC2/n218 ), .B(pgadrovfh), .C(\SAEXE/SRC2/n220 ), .D(
        \SAEXE/SRC2/n211 ) );
    snl_muxi21x1 \SAEXE/SRC2/U140  ( .ZN(\SAEXE/SRC2/n210 ), .A(
        \SAEXE/stage_1st ), .B(\SAEXE/SRC2/n208 ), .S(\SAEXE/SRC2/eqst[1] ) );
    snl_nor02x1 \SAEXE/SRC2/U100  ( .ZN(\SAEXE/srcrd_st ), .A(pgadrovfh), .B(
        \SAEXE/SRC2/n202 ) );
    snl_invx05 \SAEXE/SRC2/U112  ( .ZN(\SAEXE/SRC2/n198 ), .A(\SAEXE/seq_end )
         );
    snl_oai012x1 \SAEXE/SRC2/U135  ( .ZN(\SAEXE/SRC2/n199 ), .A(
        \SAEXE/stage_2nd ), .B(\SAEXE/SRC2/n211 ), .C(\SAEXE/SRC2/n220 ) );
    snl_nor02x1 \SAEXE/SRC2/U110  ( .ZN(\SAEXE/SRC2/n214 ), .A(
        \SAEXE/SRC2/n184 ), .B(\SAEXE/ph_lber1_h ) );
    snl_nand13x1 \SAEXE/SRC2/U127  ( .ZN(\SAEXE/SRC2/n219 ), .A(
        \SAEXE/srcwrit ), .B(\SAEXE/SRC2/n215 ), .C(\SAEXE/srcread ) );
    snl_nand12x1 \SAEXE/SRC2/U137  ( .ZN(\SAEXE/SRC2/n221 ), .A(
        \SAEXE/stage_1st ), .B(\SAEXE/SRC2/eqst[2] ) );
    snl_aoi012x1 \SAEXE/SRC2/U102  ( .ZN(\SAEXE/adovflth1 ), .A(
        \SAEXE/SRC2/n202 ), .B(\SAEXE/SRC2/n205 ), .C(\SAEXE/SRC2/n188 ) );
    snl_nand02x1 \SAEXE/SRC2/U119  ( .ZN(\SAEXE/SRC2/n217 ), .A(
        \SAEXE/stage_2nd ), .B(\SAEXE/SRC2/n206 ) );
    snl_nand02x1 \SAEXE/SRC2/U125  ( .ZN(\SAEXE/SRC2/n185 ), .A(
        \SAEXE/SRC2/n214 ), .B(\SAEXE/SRC2/n215 ) );
    snl_nor02x1 \SAEXE/SRC2/U104  ( .ZN(\SAEXE/SRC2/n207 ), .A(
        \SAEXE/SRC2/n198 ), .B(\SAEXE/SRC2/n200 ) );
    snl_aoi0b13x0 \SAEXE/SRC2/U105  ( .ZN(\SAEXE/SRC2/n187 ), .A(ph_saexe_sth), 
        .B(\SAEXE/SRC2/n208 ), .C(\SAEXE/SRC2/n209 ), .D(\SAEXE/SRC2/n210 ) );
    snl_nand13x1 \SAEXE/SRC2/U117  ( .ZN(\SAEXE/SRC2/n204 ), .A(
        \SAEXE/SRC2/eqst[4] ), .B(\SAEXE/SRC2/n213 ), .C(\SAEXE/stage_2nd ) );
    snl_oa112x1 \SAEXE/SRC2/U122  ( .Z(\SAEXE/SRC2/n189 ), .A(
        \SAEXE/ph_lber1_h ), .B(\SAEXE/SRC2/n217 ), .C(\SAEXE/SRC2/n193 ), .D(
        \SAEXE/SRC2/n218 ) );
    snl_nand02x1 \SAEXE/SRC2/U139  ( .ZN(\SAEXE/SRC2/n205 ), .A(
        \SAEXE/stage_2nd ), .B(\SAEXE/SRC2/n213 ) );
    snl_aoib122x0 \SAEXE/SRC2/U130  ( .ZN(\SAEXE/SRC2/n191 ), .A(
        \SAEXE/SRC2/n214 ), .B(\SAEXE/singlen ), .C(\SAEXE/SRC2/eqst[1] ), .D(
        \SAEXE/SRC2/n221 ), .E(\SAEXE/SRC2/n185 ) );
    snl_oai012x1 \SAEXE/SRC2/U138  ( .ZN(\SAEXE/SRC2/n222 ), .A(
        \SAEXE/SRC2/eqst[1] ), .B(\SAEXE/SRC2/n192 ), .C(\SAEXE/SRC2/n210 ) );
    snl_ffqrnx1 \SAEXE/SRC2/eqst_reg[2]  ( .Q(\SAEXE/SRC2/eqst[2] ), .D(
        \SAEXE/SRC2/nqst[2] ), .RN(n10735), .CP(SCLK) );
    snl_invx05 \SAEXE/SRC2/U116  ( .ZN(\SAEXE/SRC2/n208 ), .A(
        \SAEXE/stage_2nd ) );
    snl_nand02x1 \SAEXE/SRC2/U123  ( .ZN(\SAEXE/SRC2/n186 ), .A(
        \SAEXE/stage_1st ), .B(\SAEXE/SRC2/n206 ) );
    snl_aoi023x0 \SAEXE/SRC2/U131  ( .ZN(\SAEXE/SRC2/n190 ), .A(
        \SAEXE/SRC2/n214 ), .B(\SAEXE/singlen ), .C(\SAEXE/seq_end ), .D(
        \SAEXE/SRC2/n222 ), .E(\SAEXE/SRC2/n195 ) );
    snl_ffqrnx1 \SAEXE/SRC2/eqst_reg[4]  ( .Q(\SAEXE/SRC2/eqst[4] ), .D(
        ph_lblockh), .RN(n10735), .CP(SCLK) );
    snl_aoi1b12x0 \SAEXE/SRC2/U103  ( .ZN(\SAEXE/SRC2/n201 ), .A(
        \SAEXE/stage_2nd ), .B(\SAEXE/SRC2/n206 ), .C(\SAEXE/SRC2/n184 ), .D(
        \SAEXE/SRC2/n197 ) );
    snl_invx05 \SAEXE/SRC2/U111  ( .ZN(\SAEXE/SRC2/n215 ), .A(\SAEXE/sequen )
         );
    snl_nor02x1 \SAEXE/SRC2/U136  ( .ZN(\SAEXE/SRC2/n192 ), .A(
        \SAEXE/stage_2nd ), .B(\SAEXE/SRC2/eqst[4] ) );
    snl_invx05 \SAEXE/SRC2/U124  ( .ZN(\SAEXE/SRC2/n188 ), .A(pgadrovfh) );
    snl_invx05 \SAEXE/SRC2/U118  ( .ZN(\SAEXE/SRC2/n200 ), .A(
        \SAEXE/ph_lber1_h ) );
    snl_ffqrnx1 \SAEXE/SRC2/eqst_reg[0]  ( .Q(\SAEXE/stage_1st ), .D(
        \SAEXE/SRC2/nqst[0] ), .RN(n10735), .CP(SCLK) );
    snl_nand14x0 \MCD/rd_wt_2/U88  ( .ZN(saenabl2), .A(rrmw2), .B(
        \MCD/rd_wt_2/n4367 ), .C(\MCD/rd_wt_2/n4368 ), .D(\MCD/rd_wt_2/n4369 )
         );
    snl_ao023x1 \MCD/rd_wt_2/U89  ( .Z(ronly2), .A(\stream2[27] ), .B(
        \stream2[26] ), .C(\MCD/rd_wt_2/n4370 ), .D(\MCD/rd_wt_2/n4371 ), .E(
        \MCD/rd_wt_2/n4372 ) );
    snl_and02x1 \MCD/rd_wt_2/U90  ( .Z(po_shelter_h2), .A(\MCD/rd_wt_2/n4373 ), 
        .B(\stream2[25] ) );
    snl_aoi012x1 \MCD/rd_wt_2/U91  ( .ZN(\MCD/rd_wt_2/n4374 ), .A(
        \MCD/rd_wt_2/bacc ), .B(\stream2[1] ), .C(\MCD/rd_wt_2/n4375 ) );
    snl_nor02x1 \MCD/rd_wt_2/U96  ( .ZN(\MCD/rd_wt_2/n4373 ), .A(\stream2[27] 
        ), .B(\stream2[26] ) );
    snl_oai012x1 \MCD/rd_wt_2/U113  ( .ZN(\MCD/rd_wt_2/n4399 ), .A(
        \MCD/rd_wt_2/n4378 ), .B(\MCD/rd_wt_2/n4386 ), .C(\MCD/rd_wt_2/n4400 )
         );
    snl_invx05 \MCD/rd_wt_2/U134  ( .ZN(\MCD/rd_wt_2/n4406 ), .A(
        \MCD/rd_wt_2/n4390 ) );
    snl_invx05 \MCD/rd_wt_2/U98  ( .ZN(\MCD/rd_wt_2/n4387 ), .A(\stream2[26] )
         );
    snl_nor02x1 \MCD/rd_wt_2/U101  ( .ZN(\MCD/rd_wt_2/n4388 ), .A(
        \MCD/rd_wt_2/n4375 ), .B(\stream2[1] ) );
    snl_nand03x0 \MCD/rd_wt_2/U108  ( .ZN(\MCD/rd_wt_2/n4379 ), .A(
        \MCD/rd_wt_2/n4373 ), .B(\MCD/rd_wt_2/n4393 ), .C(\stream2[14] ) );
    snl_nor03x0 \MCD/rd_wt_2/U141  ( .ZN(\MCD/rd_wt_2/n4377 ), .A(
        \MCD/rd_wt_2/n4406 ), .B(\stream2[0] ), .C(\MCD/rd_wt_2/n4392 ) );
    snl_ffqrnx1 \MCD/rd_wt_2/ciff_reg  ( .Q(\MCD/rd_wt_2/ciff ), .D(pk_ciffh), 
        .RN(n10733), .CP(SCLK) );
    snl_nand03x0 \MCD/rd_wt_2/U106  ( .ZN(\MCD/rd_wt_2/n4392 ), .A(
        \stream2[1] ), .B(\MCD/rd_wt_2/n4375 ), .C(\MCD/rd_wt_2/n4381 ) );
    snl_and23x0 \MCD/rd_wt_2/U121  ( .Z(\MCD/rd_wt_2/n4411 ), .A(
        \MCD/rd_wt_2/n4386 ), .B(\stream2[10] ), .C(\MCD/rd_wt_2/n4373 ) );
    snl_nor02x1 \MCD/rd_wt_2/U126  ( .ZN(\MCD/rd_wt_2/n4368 ), .A(ronly2), .B(
        wonly2) );
    snl_nand14x0 \MCD/rd_wt_2/U128  ( .ZN(\MCD/rd_wt_2/n4369 ), .A(
        \stream2[22] ), .B(\MCD/rd_wt_2/n4385 ), .C(\MCD/rd_wt_2/n4372 ), .D(
        \MCD/rd_wt_2/n4399 ) );
    snl_invx05 \MCD/rd_wt_2/U146  ( .ZN(\MCD/rd_wt_2/n4402 ), .A(\stream2[18] 
        ) );
    snl_invx05 \MCD/rd_wt_2/U99  ( .ZN(\MCD/rd_wt_2/n4383 ), .A(
        \MCD/rd_wt_2/bacc ) );
    snl_aoi022x1 \MCD/rd_wt_2/U114  ( .ZN(\MCD/rd_wt_2/n4401 ), .A(
        \MCD/rd_wt_2/n4383 ), .B(\MCD/rd_wt_2/n4402 ), .C(\MCD/rd_wt_2/bacc ), 
        .D(\stream2[18] ) );
    snl_invx05 \MCD/rd_wt_2/U133  ( .ZN(sequencial2), .A(\MCD/rd_wt_2/n4392 )
         );
    snl_invx05 \MCD/rd_wt_2/U107  ( .ZN(\MCD/rd_wt_2/n4393 ), .A(\stream2[15] 
        ) );
    snl_nand02x1 \MCD/rd_wt_2/U120  ( .ZN(\MCD/rd_wt_2/n4409 ), .A(
        \MCD/rd_wt_2/n4392 ), .B(\MCD/rd_wt_2/n4410 ) );
    snl_muxi21x1 \MCD/rd_wt_2/U115  ( .ZN(\MCD/rd_wt_2/n4403 ), .A(
        \MCD/rd_wt_2/n4384 ), .B(\MCD/rd_wt_2/n4374 ), .S(\MCD/rd_wt_2/ciff )
         );
    snl_nor02x1 \MCD/rd_wt_2/U132  ( .ZN(rrmw2), .A(\MCD/rd_wt_2/n4398 ), .B(
        \MCD/rd_wt_2/n4371 ) );
    snl_xor2x0 \MCD/rd_wt_2/U95  ( .Z(\MCD/rd_wt_2/n4385 ), .A(\stream2[21] ), 
        .B(\stream2[20] ) );
    snl_invx05 \MCD/rd_wt_2/U97  ( .ZN(\MCD/rd_wt_2/n4386 ), .A(\stream2[9] )
         );
    snl_invx05 \MCD/rd_wt_2/U109  ( .ZN(\MCD/rd_wt_2/n4394 ), .A(\stream2[13] 
        ) );
    snl_invx05 \MCD/rd_wt_2/U129  ( .ZN(rmw12), .A(\MCD/rd_wt_2/n4369 ) );
    snl_invx05 \MCD/rd_wt_2/U140  ( .ZN(\MCD/rd_wt_2/n4371 ), .A(
        \MCD/rd_wt_2/n4399 ) );
    snl_invx05 \MCD/rd_wt_2/U100  ( .ZN(\MCD/rd_wt_2/n4375 ), .A(\stream2[2] )
         );
    snl_oai113x0 \MCD/rd_wt_2/U112  ( .ZN(\MCD/rd_wt_2/n4398 ), .A(
        \MCD/rd_wt_2/n4390 ), .B(\stream2[0] ), .C(\MCD/rd_wt_2/n4380 ), .D(
        \MCD/rd_wt_2/n4372 ), .E(\MCD/rd_wt_2/n4397 ) );
    snl_invx05 \MCD/rd_wt_2/U135  ( .ZN(\MCD/rd_wt_2/n4384 ), .A(
        \MCD/rd_wt_2/n4388 ) );
    snl_oai013x0 \MCD/rd_wt_2/U110  ( .ZN(\MCD/rd_wt_2/n4372 ), .A(
        \MCD/rd_wt_2/n4393 ), .B(\MCD/rd_wt_2/n4395 ), .C(\MCD/rd_wt_2/n4377 ), 
        .D(\MCD/rd_wt_2/n4396 ) );
    snl_and34x0 \MCD/rd_wt_2/U127  ( .Z(wonly2), .A(\MCD/rd_wt_2/n4372 ), .B(
        \MCD/rd_wt_2/n4371 ), .C(\stream2[22] ), .D(\MCD/rd_wt_2/n4385 ) );
    snl_invx05 \MCD/rd_wt_2/U137  ( .ZN(\MCD/rd_wt_2/n4395 ), .A(
        \MCD/rd_wt_2/n4409 ) );
    snl_invx05 \MCD/rd_wt_2/U102  ( .ZN(\MCD/rd_wt_2/n4389 ), .A(\stream2[0] )
         );
    snl_aoi222x0 \MCD/rd_wt_2/U119  ( .ZN(\MCD/rd_wt_2/n4408 ), .A(
        \MCD/rd_wt_2/n4375 ), .B(\MCD/rd_wt_2/n4391 ), .C(\MCD/rd_wt_2/n4388 ), 
        .D(\MCD/rd_wt_2/n4383 ), .E(\stream2[1] ), .F(\MCD/rd_wt_2/n4390 ) );
    snl_aoi022x1 \MCD/rd_wt_2/U142  ( .ZN(\MCD/rd_wt_2/n4415 ), .A(
        \MCD/rd_wt_2/n4405 ), .B(\MCD/rd_wt_2/n4389 ), .C(\MCD/rd_wt_2/n4404 ), 
        .D(\stream2[0] ) );
    snl_aoi012x1 \MCD/rd_wt_2/U125  ( .ZN(\MCD/rd_wt_2/n4370 ), .A(
        \stream2[19] ), .B(\MCD/rd_wt_2/n4401 ), .C(\stream2[25] ) );
    snl_nor02x1 \MCD/rd_wt_2/U105  ( .ZN(\MCD/rd_wt_2/n4381 ), .A(
        \MCD/rd_wt_2/n4387 ), .B(\stream2[27] ) );
    snl_nor02x1 \MCD/rd_wt_2/U122  ( .ZN(\MCD/rd_wt_2/n4412 ), .A(
        \stream2[13] ), .B(\MCD/rd_wt_2/n4379 ) );
    snl_oa113x1 \MCD/rd_wt_2/U139  ( .Z(\MCD/rd_wt_2/n4378 ), .A(
        \MCD/rd_wt_2/n4414 ), .B(\MCD/rd_wt_2/n4380 ), .C(\MCD/rd_wt_2/n4389 ), 
        .D(\MCD/rd_wt_2/n4392 ), .E(\MCD/rd_wt_2/n4416 ) );
    snl_oa012x1 \MCD/rd_wt_2/U92  ( .Z(\MCD/rd_wt_2/n4376 ), .A(
        \MCD/rd_wt_2/n4377 ), .B(\MCD/rd_wt_2/n4378 ), .C(\MCD/rd_wt_2/n4379 )
         );
    snl_muxi21x1 \MCD/rd_wt_2/U145  ( .ZN(\MCD/rd_wt_2/n4396 ), .A(
        \MCD/rd_wt_2/n4413 ), .B(\MCD/rd_wt_2/n4412 ), .S(\stream2[12] ) );
    snl_nand02x1 \MCD/rd_wt_2/U93  ( .ZN(\MCD/rd_wt_2/n4380 ), .A(
        \MCD/rd_wt_2/n4381 ), .B(\stream2[1] ) );
    snl_invx05 \MCD/rd_wt_2/U104  ( .ZN(\MCD/rd_wt_2/n4391 ), .A(pk_sign_h) );
    snl_aoi222x0 \MCD/rd_wt_2/U117  ( .ZN(\MCD/rd_wt_2/n4405 ), .A(pk_sign_h), 
        .B(\MCD/rd_wt_2/n4375 ), .C(\MCD/rd_wt_2/n4388 ), .D(
        \MCD/rd_wt_2/bacc ), .E(\MCD/rd_wt_2/n4406 ), .F(\stream2[1] ) );
    snl_nand03x0 \MCD/rd_wt_2/U130  ( .ZN(\MCD/rd_wt_2/n4367 ), .A(
        \MCD/rd_wt_2/n4398 ), .B(\MCD/rd_wt_2/n4399 ), .C(\MCD/rd_wt_2/n4397 )
         );
    snl_nand02x1 \MCD/rd_wt_2/U138  ( .ZN(\MCD/rd_wt_2/n4416 ), .A(
        \MCD/rd_wt_2/n4417 ), .B(\MCD/rd_wt_2/n4381 ) );
    snl_aoi013x0 \MCD/rd_wt_2/U116  ( .ZN(\MCD/rd_wt_2/n4404 ), .A(ph_piosl_h), 
        .B(\pk_stat_h[18] ), .C(\stream2[1] ), .D(\MCD/rd_wt_2/n4403 ) );
    snl_nor02x1 \MCD/rd_wt_2/U123  ( .ZN(\MCD/rd_wt_2/n4413 ), .A(
        \MCD/rd_wt_2/n4376 ), .B(\MCD/rd_wt_2/n4394 ) );
    snl_invx05 \MCD/rd_wt_2/U131  ( .ZN(rmw22), .A(\MCD/rd_wt_2/n4367 ) );
    snl_ffqrnx1 \MCD/rd_wt_2/bacc_reg  ( .Q(\MCD/rd_wt_2/bacc ), .D(pk_bacch), 
        .RN(n10733), .CP(SCLK) );
    snl_nor02x1 \MCD/rd_wt_2/U94  ( .ZN(\MCD/rd_wt_2/n4382 ), .A(
        \MCD/rd_wt_2/n4383 ), .B(\MCD/rd_wt_2/n4384 ) );
    snl_aoi022x1 \MCD/rd_wt_2/U143  ( .ZN(\MCD/rd_wt_2/n4417 ), .A(
        \MCD/rd_wt_2/n4408 ), .B(\MCD/rd_wt_2/n4389 ), .C(\MCD/rd_wt_2/n4407 ), 
        .D(\stream2[0] ) );
    snl_muxi21x1 \MCD/rd_wt_2/U144  ( .ZN(\MCD/rd_wt_2/n4400 ), .A(
        \MCD/rd_wt_2/n4411 ), .B(\MCD/rd_wt_2/n4409 ), .S(\stream2[11] ) );
    snl_nand12x1 \MCD/rd_wt_2/U103  ( .ZN(\MCD/rd_wt_2/n4390 ), .A(pk_pcon31_h
        ), .B(\MCD/rd_wt_2/ciff ) );
    snl_nor03x0 \MCD/rd_wt_2/U111  ( .ZN(\MCD/rd_wt_2/n4397 ), .A(
        \stream2[22] ), .B(\stream2[20] ), .C(\stream2[21] ) );
    snl_nand02x1 \MCD/rd_wt_2/U136  ( .ZN(\MCD/rd_wt_2/n4410 ), .A(
        \MCD/rd_wt_2/n4415 ), .B(\MCD/rd_wt_2/n4381 ) );
    snl_ao022x1 \MCD/rd_wt_2/U124  ( .Z(\MCD/rd_wt_2/n4414 ), .A(
        \MCD/rd_wt_2/bacc ), .B(\MCD/rd_wt_2/ciff ), .C(\pk_stat_h[18] ), .D(
        ph_piosl_h) );
    snl_muxi21x1 \MCD/rd_wt_2/U118  ( .ZN(\MCD/rd_wt_2/n4407 ), .A(
        \MCD/rd_wt_2/n4375 ), .B(\MCD/rd_wt_2/n4382 ), .S(\MCD/rd_wt_2/ciff )
         );
    snl_invx2 \REGF/pbmemff41/U1225  ( .ZN(\REGF/pbmemff41/n7083 ), .A(
        \REGF/pbmemff41/n7082 ) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[20]  ( .Q(CDOUT[52]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOH[20] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[13]  ( .Q(CDOUT[45]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\REGF/RI_PCOH[13] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[5]  ( .Q(\REGF/RO_SRDA[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRDA[5] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[1]  ( .Q(\pk_sra2_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[1] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[20]  ( .Q(\pk_s01l_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[13]  ( .Q(\pk_s01l_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[26]  ( .Q(\pk_sefl_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[15]  ( .Q(\pk_sefl_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[6]  ( .Q(\pk_s23l_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[31]  ( .Q(\pk_sabl_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[28]  ( .Q(\pk_sabl_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[21]  ( .Q(\pk_s23l_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[12]  ( .Q(\pk_s23l_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1242  ( .ZN(\REGF/pbmemff41/n7099 ), .A(
        \REGF/pbmemff41/n7097 ) );
    snl_and02x1 \REGF/pbmemff41/U1250  ( .Z(\REGF/pbmemff41/RO_PSAS9B551[4] ), 
        .A(ph_lbe3_h), .B(\REGF/pbmemff41/n7103 ) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[5]  ( .Q(CDOUT[37]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOH[5] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[19]  ( .Q(\pk_s89l_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[8]  ( .Q(\pk_sra2_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[8] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[6]  ( .Q(\pk_s01l_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[31]  ( .Q(\pk_s23l_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[26]  ( .Q(\pk_s67l_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[15]  ( .Q(\pk_s67l_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[6]  ( .Q(\pk_sefl_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[28]  ( .Q(\pk_s23l_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[20]  ( .Q(\REGF/RO_ERRA[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\pgsadrh[20] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[10]  ( .Q(\pk_s89l_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[13]  ( .Q(\REGF/RO_ERRA[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\pgsadrh[13] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[23]  ( .Q(\pk_s89l_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[6]  ( .Q(\pk_trba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_TBAI[6] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[30]  ( .Q(\pk_s01l_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[21]  ( .Q(\pk_sabl_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[29]  ( .Q(\pk_s01l_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[12]  ( .Q(\pk_sabl_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1277  ( .Z(
        \REGF/pbmemff41/*cell*5493/U16/DATA2_0 ), .A(PDLIN[4]), .B(\pgldi[4] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[27]  ( .Q(\pk_s45l_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[1]  ( .Q(CDOUT[33]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\REGF/RI_PCOH[1] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[14]  ( .Q(\pk_s45l_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1265  ( .Z(
        \REGF/pbmemff41/*cell*5493/U67/Z_0 ), .A(PDLIN[23]), .B(\pgldi[7] ), 
        .S(ph_tbllt_h) );
    snl_mux21x1 \REGF/pbmemff41/U1280  ( .Z(
        \REGF/pbmemff41/*cell*5493/U10/DATA2_0 ), .A(PDLIN[7]), .B(\pgldi[7] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[5]  ( .Q(\pk_sra2_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_SRA12M[5] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[16]  ( .Q(\pk_s23l_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[18]  ( .Q(\pk_s67l_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[25]  ( .Q(\pk_s23l_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[24]  ( .Q(\pk_s01l_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[17]  ( .Q(\pk_s01l_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[2]  ( .Q(\pk_s23l_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[19]  ( .Q(\pk_s45l_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[11]  ( .Q(\pk_sefl_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_bufx1 \REGF/pbmemff41/U1224  ( .Z(\REGF/pbmemff41/n7082 ), .A(
        \REGF/pbmemff41/n7102 ) );
    snl_invx2 \REGF/pbmemff41/U1230  ( .ZN(\REGF/pbmemff41/n7088 ), .A(
        \REGF/pbmemff41/n7087 ) );
    snl_invx2 \REGF/pbmemff41/U1237  ( .ZN(\REGF/pbmemff41/n7094 ), .A(
        \REGF/pbmemff41/n7092 ) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[24]  ( .Q(CDOUT[56]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[24] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[1]  ( .Q(\REGF/RO_SRDA[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRDA[1] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[22]  ( .Q(\pk_sefl_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[17]  ( .Q(CDOUT[49]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOH[17] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1259  ( .Z(
        \REGF/pbmemff41/*cell*5493/U79/Z_0 ), .A(PDLIN[17]), .B(\pgldi[1] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[8]  ( .Q(CDOUT[40]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[8] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[8]  ( .Q(\REGF/RO_SRDA[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRDA[8] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[2]  ( .Q(\pk_trba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_TBAI[2] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[23]  ( .Q(\pk_s45l_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[10]  ( .Q(\pk_s45l_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[25]  ( .Q(\pk_sabl_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[18]  ( .Q(\pk_sefl_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[16]  ( .Q(\pk_sabl_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[24]  ( .Q(\REGF/RO_ERRA[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\pgsadrh[24] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[17]  ( .Q(\REGF/RO_ERRA[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\pgsadrh[17] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[14]  ( .Q(\pk_s89l_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[27]  ( .Q(\pk_s89l_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[2]  ( .Q(\pk_sefl_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1279  ( .Z(
        \REGF/pbmemff41/*cell*5493/U12/DATA2_0 ), .A(PDLIN[6]), .B(\pgldi[6] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[26]  ( .Q(\REGF/RO_ERRA[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\pgsadrh[26] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[2]  ( .Q(\pk_s01l_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[22]  ( .Q(\pk_s67l_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[11]  ( .Q(\pk_s67l_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[16]  ( .Q(\pk_s89l_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[15]  ( .Q(\REGF/RO_ERRA[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[15] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[25]  ( .Q(\pk_s89l_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[0]  ( .Q(\pk_s01l_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[20]  ( .Q(\pk_s67l_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[9]  ( .Q(\pk_s23l_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[21]  ( .Q(\pk_s45l_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[13]  ( .Q(\pk_s67l_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[0]  ( .Q(\pk_sefl_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[12]  ( .Q(\pk_s45l_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[30]  ( .Q(\pk_sefl_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[29]  ( .Q(\pk_sefl_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[27]  ( .Q(\pk_sabl_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[14]  ( .Q(\pk_sabl_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1231  ( .ZN(\REGF/pbmemff41/n7091 ), .A(
        \REGF/pbmemff41/n7087 ) );
    snl_bufx1 \REGF/pbmemff41/U1239  ( .Z(\REGF/pbmemff41/n7097 ), .A(
        \REGF/pbmemff41/n7102 ) );
    snl_or02x1 \REGF/pbmemff41/U1245  ( .Z(
        \REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), .A(ph_tpralt_h), .B(
        \pk_rwrit_h[46] ) );
    snl_mux21x1 \REGF/pbmemff41/U1262  ( .Z(
        \REGF/pbmemff41/*cell*5493/U73/Z_0 ), .A(PDLIN[20]), .B(\pgldi[4] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[26]  ( .Q(CDOUT[58]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOH[26] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[0]  ( .Q(\pk_trba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_TBAI[0] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[26]  ( .Q(\pk_s01l_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[15]  ( .Q(\pk_s01l_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[0]  ( .Q(\pk_s23l_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[31]  ( .Q(\pk_s45l_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[28]  ( .Q(\pk_s45l_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[13]  ( .Q(\pk_sefl_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[20]  ( .Q(\pk_sefl_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[15]  ( .Q(CDOUT[47]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[15] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[3]  ( .Q(\REGF/RO_SRDA[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[3] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[9]  ( .Q(\pk_trba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_TBAI[9] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[3]  ( .Q(CDOUT[35]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOH[3] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1257  ( .Z(
        \REGF/pbmemff41/*cell*5493/U81/Z_0 ), .A(PDLIN[16]), .B(\pgldi[0] ), 
        .S(ph_tbllt_h) );
    snl_mux21x1 \REGF/pbmemff41/U1270  ( .Z(
        \REGF/pbmemff41/*cell*5493/U59/Z_0 ), .A(PDLIN[27]), .B(\pgldi[11] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[18]  ( .Q(CDOUT[50]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOH[18] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[7]  ( .Q(\pk_sra2_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[7] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[9]  ( .Q(\pk_s01l_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[30]  ( .Q(\pk_s67l_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[29]  ( .Q(\pk_s67l_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[9]  ( .Q(\pk_sefl_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[27]  ( .Q(\pk_s23l_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[14]  ( .Q(\pk_s23l_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[4]  ( .Q(\pk_trba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_TBAI[4] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[23]  ( .Q(\pk_sabl_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[18]  ( .Q(\pk_s01l_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[10]  ( .Q(\pk_sabl_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[25]  ( .Q(\pk_s45l_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[16]  ( .Q(\pk_s45l_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[4]  ( .Q(\pk_sefl_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_invx1 \REGF/pbmemff41/U1244  ( .ZN(\REGF/pbmemff41/n7102 ), .A(
        \REGF/n8052 ) );
    snl_mux21x1 \REGF/pbmemff41/U1263  ( .Z(
        \REGF/pbmemff41/*cell*5493/U71/Z_0 ), .A(PDLIN[21]), .B(\pgldi[5] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[22]  ( .Q(CDOUT[54]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOH[22] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[7]  ( .Q(CDOUT[39]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[7] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[3]  ( .Q(\pk_sra2_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[3] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[22]  ( .Q(\REGF/RO_ERRA[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[22] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[4]  ( .Q(\pk_s01l_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[24]  ( .Q(\pk_s67l_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[19]  ( .Q(\pk_s23l_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[17]  ( .Q(\pk_s67l_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[11]  ( .Q(\REGF/RO_ERRA[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\pgsadrh[11] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[12]  ( .Q(\pk_s89l_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[10]  ( .Q(\pk_s23l_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[21]  ( .Q(\pk_s89l_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[18]  ( .Q(\REGF/RO_ERRA[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\pgsadrh[18] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[23]  ( .Q(\pk_s23l_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[31]  ( .Q(\pk_s89l_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[28]  ( .Q(\pk_s89l_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[7]  ( .Q(\REGF/RO_SRDA[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[7] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[11]  ( .Q(CDOUT[43]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOH[11] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[4]  ( .Q(\pk_sra1_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRA12M[4] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[22]  ( .Q(\pk_s01l_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[11]  ( .Q(\pk_s01l_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[19]  ( .Q(\pk_sabl_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[24]  ( .Q(\pk_sefl_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[17]  ( .Q(\pk_sefl_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[4]  ( .Q(\pk_s23l_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[5]  ( .Q(\pk_s89l_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[23]  ( .Q(CDOUT[23]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[23] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[19]  ( .Q(CDOUT[19]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOL[19] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[22]  ( .Q(\pk_sra1_h[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[22] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[4]  ( .Q(\pk_s45l_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[4]  ( .Q(\pk_sabl_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[11]  ( .Q(\pk_sra1_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_SRA12M[11] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[26]  ( .Q(\pk_sra2_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[26] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[26]  ( .Q(\REGF/RO_SRDA[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRDA[26] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[0]  ( .Q(\pk_scdl_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[10]  ( .Q(CDOUT[10]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[10] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[3]  ( .Q(CDOUT[3]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[3] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[15]  ( .Q(\pk_sra2_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[15] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[15]  ( .Q(\REGF/RO_SRDA[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_SRDA[15] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[5]  ( .Q(\REGF/RO_EST1[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(
        \REGF/pbmemff41/RO_PSAS9B551[5] ), .SE(\REGF/pbmemff41/n_2861 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[14]  ( .Q(\pk_stdat[14] ), .D(
        \REGF/pbmemff41/*cell*5493/U77/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7091 ), .SD(\REGF/pbmemff41/RO_TRCOT[14] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[7]  ( .Q(\pk_stdat[7] ), .D(
        \REGF/pbmemff41/*cell*5493/U10/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7098 ), .SD(\REGF/pbmemff41/RO_TRCOT[7] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1238  ( .ZN(\REGF/pbmemff41/n7095 ), .A(
        \REGF/pbmemff41/n7092 ) );
    snl_mux21x1 \REGF/pbmemff41/U1278  ( .Z(
        \REGF/pbmemff41/*cell*5493/U14/DATA2_0 ), .A(PDLIN[5]), .B(\pgldi[5] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[18]  ( .Q(\pk_sra1_h[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[18] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[1]  ( .Q(\pk_psae_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[4]  ( .Q(\pk_s67l_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[9]  ( .Q(\pk_scdl_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[5]  ( .Q(\REGF/RO_ERRA[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[5] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[15]  ( .Q(\pk_scdl_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[17]  ( .Q(\pk_trba_h[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_TBAI[17] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[26]  ( .Q(\pk_scdl_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[7]  ( .Q(CDOUT[7]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[7] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[22]  ( .Q(\pk_sra2_h[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[22] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[9]  ( .Q(\pk_s67l_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[8]  ( .Q(\REGF/RO_PSASH[15] ), 
        .D(ph_trsc_h), .EN(\REGF/pbmemff41/n8037 ), .RN(\REGF/pbmemff41/n7090 
        ), .SD(1'b0), .SE(\pk_rwrit_h[48] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[19]  ( .Q(\pk_stdat[19] ), .D(
        \REGF/pbmemff41/*cell*5493/U67/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7100 ), .SD(\REGF/pbmemff41/RO_TRCOT[19] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[22]  ( .Q(\REGF/RO_SRDA[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRDA[22] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[4]  ( .Q(\pk_scdl_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[26]  ( .Q(\pk_sra1_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[26] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[11]  ( .Q(\pk_sra2_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[11] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[11]  ( .Q(\REGF/RO_SRDA[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[11] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[15]  ( .Q(\pk_sra1_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[15] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[0]  ( .Q(\pk_sra1_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_SRA12M[0] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[8]  ( .Q(\REGF/RO_ERRA[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\pgsadrh[8] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[18]  ( .Q(\pk_scdl_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[0]  ( .Q(\pk_s45l_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[0]  ( .Q(\pk_sabl_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[1]  ( .Q(\pk_s89l_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_nand12x1 \REGF/pbmemff41/U1251  ( .ZN(\REGF/pbmemff41/n_2859 ), .A(
        phsaerrh), .B(\REGF/pbmemff41/n7103 ) );
    snl_nor02x1 \REGF/pbmemff41/U1256  ( .ZN(\REGF/pbmemff41/n7103 ), .A(
        \pk_rwrit_h[48] ), .B(\pk_rwrit_h[55] ) );
    snl_mux21x1 \REGF/pbmemff41/U1271  ( .Z(
        \REGF/pbmemff41/*cell*5493/U4/DATA2_0 ), .A(PDLIN[10]), .B(\pgldi[10] 
        ), .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[14]  ( .Q(CDOUT[14]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOL[14] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[9]  ( .Q(\pk_sra1_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[9] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[1]  ( .Q(\REGF/RO_ERRA[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[1] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[20]  ( .Q(\pk_trba_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_TBAI[20] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[13]  ( .Q(\pk_trba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_TBAI[13] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[11]  ( .Q(\pk_scdl_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[8]  ( .Q(\pk_s89l_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[22]  ( .Q(\pk_scdl_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[18]  ( .Q(\pk_sra2_h[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[18] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[5]  ( .Q(\pk_psae_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[9]  ( .Q(\pk_s45l_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[9]  ( .Q(\pk_sabl_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[0]  ( .Q(\pk_s67l_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[18]  ( .Q(\REGF/RO_SRDA[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[18] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[27]  ( .Q(CDOUT[27]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOL[27] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[23]  ( .Q(\REGF/RO_TRCO[27] ), 
        .D(\REGF/pbmemff41/*cell*5493/U59/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7099 ), .SD(\REGF/pbmemff41/RO_TRCOT[23] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[25]  ( .Q(CDOUT[25]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOL[25] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[16]  ( .Q(CDOUT[16]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOL[16] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[2]  ( .Q(\pk_s67l_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[1]  ( .Q(\REGF/RO_PSASL[1] ), 
        .D(ph_tcer_h), .EN(\REGF/pbmemff41/n8037 ), .RN(\REGF/pbmemff41/n7090 
        ), .SD(1'b0), .SE(\pk_rwrit_h[48] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[10]  ( .Q(\pk_stdat[10] ), .D(
        \REGF/pbmemff41/*cell*5493/U4/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7090 ), .SD(\REGF/pbmemff41/RO_TRCOT[10] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[3]  ( .Q(\pk_stdat[3] ), .D(
        \REGF/pbmemff41/*cell*5493/U18/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7098 ), .SD(\REGF/pbmemff41/RO_TRCOT[3] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1276  ( .Z(
        \REGF/pbmemff41/*cell*5493/U18/DATA2_0 ), .A(PDLIN[3]), .B(\pgldi[3] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[30]  ( .Q(\REGF/RO_SRDA[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_SRDA[30] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[29]  ( .Q(\REGF/RO_SRDA[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRDA[29] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[3]  ( .Q(\REGF/RO_EST1[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(
        \REGF/pbmemff41/RO_PSAS9B551[3] ), .SE(\REGF/pbmemff41/n_2859 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[24]  ( .Q(\pk_sra1_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[24] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[7]  ( .Q(\pk_psae_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[3]  ( .Q(\REGF/RO_ERRA[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\pgsadrh[3] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[13]  ( .Q(\pk_scdl_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[21]  ( .Q(\REGF/RO_TRCO[25] ), 
        .D(\REGF/pbmemff41/*cell*5493/U63/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7099 ), .SD(\REGF/pbmemff41/RO_TRCOT[21] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[12]  ( .Q(\pk_stdat[12] ), .D(
        \REGF/pbmemff41/*cell*5493/U81/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7088 ), .SD(\REGF/pbmemff41/RO_TRCOT[12] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[1]  ( .Q(\pk_stdat[1] ), .D(
        \REGF/pbmemff41/*cell*5493/U22/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7099 ), .SD(\REGF/pbmemff41/RO_TRCOT[1] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[22]  ( .Q(\pk_trba_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_TBAI[22] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[11]  ( .Q(\pk_trba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_TBAI[11] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[20]  ( .Q(\pk_scdl_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[30]  ( .Q(\pk_scdl_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[29]  ( .Q(\pk_scdl_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[17]  ( .Q(\pk_sra1_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[17] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[18]  ( .Q(\pk_trba_h[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_TBAI[18] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1226  ( .ZN(\REGF/pbmemff41/n7086 ), .A(
        \REGF/pbmemff41/n7082 ) );
    snl_invx2 \REGF/pbmemff41/U1236  ( .ZN(\REGF/pbmemff41/n7096 ), .A(
        \REGF/pbmemff41/n7092 ) );
    snl_mux21x1 \REGF/pbmemff41/U1258  ( .Z(
        \REGF/pbmemff41/*cell*5493/U8/DATA2_0 ), .A(PDLIN[8]), .B(\pgldi[8] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[5]  ( .Q(CDOUT[5]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOL[5] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[2]  ( .Q(\pk_sra1_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[2] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[2]  ( .Q(\pk_s45l_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[3]  ( .Q(\pk_s89l_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[2]  ( .Q(\pk_sabl_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[20]  ( .Q(\pk_sra2_h[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[20] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[20]  ( .Q(\REGF/RO_SRDA[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[20] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[6]  ( .Q(\pk_scdl_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[8]  ( .Q(\pk_stdat[8] ), .D(
        \REGF/pbmemff41/*cell*5493/U8/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7090 ), .SD(\REGF/pbmemff41/RO_TRCOT[8] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[13]  ( .Q(\pk_sra2_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[13] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[13]  ( .Q(\REGF/RO_SRDA[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_SRDA[13] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[3]  ( .Q(\pk_psae_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[7]  ( .Q(\REGF/RO_ERRA[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[7] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[15]  ( .Q(\pk_trba_h[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_TBAI[15] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[17]  ( .Q(\pk_scdl_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[24]  ( .Q(\pk_scdl_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[7]  ( .Q(\REGF/RO_PSASL[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(ph_bitsrc_h), 
        .SE(ad_latch), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1243  ( .ZN(\REGF/pbmemff41/n7100 ), .A(
        \REGF/pbmemff41/n7097 ) );
    snl_nor02x1 \REGF/pbmemff41/U1281  ( .ZN(\REGF/pbmemff41/n8035 ), .A(
        \pk_rwrit_h[45] ), .B(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[21]  ( .Q(CDOUT[21]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOL[21] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[12]  ( .Q(CDOUT[12]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[12] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[8]  ( .Q(CDOUT[8]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOL[8] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[16]  ( .Q(\pk_stdat[16] ), .D(
        \REGF/pbmemff41/*cell*5493/U73/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7090 ), .SD(\REGF/pbmemff41/RO_TRCOT[16] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[5]  ( .Q(\pk_stdat[5] ), .D(
        \REGF/pbmemff41/*cell*5493/U14/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7100 ), .SD(\REGF/pbmemff41/RO_TRCOT[5] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[24]  ( .Q(\pk_sra2_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[24] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[6]  ( .Q(\pk_s67l_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[24]  ( .Q(\REGF/RO_SRDA[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRDA[24] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[2]  ( .Q(\pk_scdl_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[31]  ( .Q(CDOUT[31]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[31] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[28]  ( .Q(CDOUT[28]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\REGF/RI_PCOL[28] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[1]  ( .Q(CDOUT[1]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\REGF/RI_PCOL[1] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[17]  ( .Q(\pk_sra2_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[17] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[17]  ( .Q(\REGF/RO_SRDA[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_SRDA[17] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_and02x1 \REGF/pbmemff41/U1248  ( .Z(\REGF/pbmemff41/RO_PSAS9B551[5] ), 
        .A(\REGF/D2_HINT ), .B(\REGF/pbmemff41/n7103 ) );
    snl_mux21x1 \REGF/pbmemff41/U1264  ( .Z(
        \REGF/pbmemff41/*cell*5493/U69/Z_0 ), .A(PDLIN[22]), .B(\pgldi[6] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[6]  ( .Q(\pk_sra1_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRA12M[6] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[7]  ( .Q(\pk_s89l_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[20]  ( .Q(\pk_sra1_h[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[20] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[6]  ( .Q(\pk_s45l_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[6]  ( .Q(\pk_sabl_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[13]  ( .Q(\pk_sra1_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[13] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[2]  ( .Q(\pk_psae_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[20]  ( .Q(CDOUT[20]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOL[20] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[13]  ( .Q(CDOUT[13]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\REGF/RI_PCOL[13] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[6]  ( .Q(\REGF/RO_ERRA[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\pgsadrh[6] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[16]  ( .Q(\pk_scdl_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[14]  ( .Q(\pk_trba_h[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_TBAI[14] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[25]  ( .Q(\pk_scdl_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[9]  ( .Q(CDOUT[9]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOL[9] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[6]  ( .Q(\REGF/RO_PSASL[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(ph_lbwrh), .SE(
        ph_sdirlth), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1241  ( .ZN(\REGF/pbmemff41/n7101 ), .A(
        \REGF/pbmemff41/n7097 ) );
    snl_and02x1 \REGF/pbmemff41/U1253  ( .Z(\REGF/pbmemff41/RO_PSAS9B551[2] ), 
        .A(ph_lbe1_h), .B(\REGF/pbmemff41/n7103 ) );
    snl_mux21x1 \REGF/pbmemff41/U1274  ( .Z(
        \REGF/pbmemff41/*cell*5493/U20/DATA2_0 ), .A(PDLIN[2]), .B(\pgldi[2] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[30]  ( .Q(CDOUT[30]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOL[30] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[7]  ( .Q(\pk_s67l_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[17]  ( .Q(\pk_stdat[17] ), .D(
        \REGF/pbmemff41/*cell*5493/U71/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7098 ), .SD(\REGF/pbmemff41/RO_TRCOT[17] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[4]  ( .Q(\pk_stdat[4] ), .D(
        \REGF/pbmemff41/*cell*5493/U16/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7089 ), .SD(\REGF/pbmemff41/RO_TRCOT[4] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[29]  ( .Q(CDOUT[29]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOL[29] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[0]  ( .Q(CDOUT[0]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOL[0] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[25]  ( .Q(\pk_sra2_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[25] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[25]  ( .Q(\REGF/RO_SRDA[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRDA[25] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[3]  ( .Q(\pk_scdl_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[16]  ( .Q(\pk_sra2_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[16] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[16]  ( .Q(\REGF/RO_SRDA[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[16] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[7]  ( .Q(\pk_s45l_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[7]  ( .Q(\pk_sabl_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1266  ( .Z(
        \REGF/pbmemff41/*cell*5493/U65/Z_0 ), .A(PDLIN[24]), .B(\pgldi[8] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[21]  ( .Q(\pk_sra1_h[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[21] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[7]  ( .Q(\pk_sra1_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_SRA12M[7] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[6]  ( .Q(\pk_s89l_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[12]  ( .Q(\pk_sra1_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[12] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[3]  ( .Q(\pk_s67l_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[2]  ( .Q(\REGF/RO_EST1[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(
        \REGF/pbmemff41/RO_PSAS9B551[2] ), .SE(\REGF/pbmemff41/n_2859 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[20]  ( .Q(\pk_stdat[20] ), .D(
        \REGF/pbmemff41/*cell*5493/U65/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7088 ), .SD(\REGF/pbmemff41/RO_TRCOT[20] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[24]  ( .Q(CDOUT[24]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOL[24] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[17]  ( .Q(CDOUT[17]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOL[17] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[13]  ( .Q(\pk_stdat[13] ), .D(
        \REGF/pbmemff41/*cell*5493/U79/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7098 ), .SD(\REGF/pbmemff41/RO_TRCOT[13] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[0]  ( .Q(\pk_stdat[0] ), .D(
        \REGF/pbmemff41/*cell*5493/U24/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7089 ), .SD(\REGF/pbmemff41/RO_TRCOT[0] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[31]  ( .Q(\REGF/RO_SRDA[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRDA[31] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[28]  ( .Q(\REGF/RO_SRDA[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRDA[28] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[6]  ( .Q(\pk_psae_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[2]  ( .Q(\REGF/RO_ERRA[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\pgsadrh[2] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[23]  ( .Q(\pk_trba_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_TBAI[23] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[10]  ( .Q(\pk_trba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_TBAI[10] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[12]  ( .Q(\pk_scdl_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[21]  ( .Q(\pk_scdl_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1227  ( .ZN(\REGF/pbmemff41/n7084 ), .A(
        \REGF/pbmemff41/n7082 ) );
    snl_invx2 \REGF/pbmemff41/U1228  ( .ZN(\REGF/pbmemff41/n7085 ), .A(
        \REGF/pbmemff41/n7082 ) );
    snl_invx2 \REGF/pbmemff41/U1233  ( .ZN(\REGF/pbmemff41/n7090 ), .A(
        \REGF/pbmemff41/n7087 ) );
    snl_bufx1 \REGF/pbmemff41/U1234  ( .Z(\REGF/pbmemff41/n7092 ), .A(
        \REGF/pbmemff41/n7102 ) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[25]  ( .Q(\pk_sra1_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[25] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[16]  ( .Q(\pk_sra1_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[16] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[19]  ( .Q(\pk_trba_h[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_TBAI[19] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[31]  ( .Q(\pk_scdl_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[28]  ( .Q(\pk_scdl_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[3]  ( .Q(\pk_sra1_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_SRA12M[3] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[2]  ( .Q(\pk_s89l_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[6]  ( .Q(CDOUT[6]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOL[6] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[4]  ( .Q(CDOUT[4]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOL[4] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[21]  ( .Q(\pk_sra2_h[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[21] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[3]  ( .Q(\pk_s45l_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[3]  ( .Q(\pk_sabl_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[7]  ( .Q(\pk_scdl_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[12]  ( .Q(\pk_sra2_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRA12M[12] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[21]  ( .Q(\REGF/RO_SRDA[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRDA[21] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[12]  ( .Q(\REGF/RO_SRDA[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_SRDA[12] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[23]  ( .Q(\pk_sra2_h[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[23] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[23]  ( .Q(\REGF/RO_SRDA[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRDA[23] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[8]  ( .Q(\pk_s67l_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[9]  ( .Q(\pk_stdat[9] ), .D(
        \REGF/pbmemff41/*cell*5493/U6/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7100 ), .SD(\REGF/pbmemff41/RO_TRCOT[9] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[5]  ( .Q(\pk_scdl_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[27]  ( .Q(\pk_sra1_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[27] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[10]  ( .Q(\pk_sra2_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[10] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[10]  ( .Q(\REGF/RO_SRDA[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[10] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[18]  ( .Q(\pk_stdat[18] ), .D(
        \REGF/pbmemff41/*cell*5493/U69/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7091 ), .SD(\REGF/pbmemff41/RO_TRCOT[18] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[14]  ( .Q(\pk_sra1_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[14] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[9]  ( .Q(\REGF/RO_ERRA[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[9] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[19]  ( .Q(\pk_scdl_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[1]  ( .Q(\pk_sra1_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[1] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[0]  ( .Q(\REGF/RO_ERRA[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[0] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[1]  ( .Q(\pk_s45l_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[0]  ( .Q(\pk_s89l_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[1]  ( .Q(\pk_sabl_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[10]  ( .Q(\pk_scdl_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[21]  ( .Q(\pk_trba_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_TBAI[21] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[12]  ( .Q(\pk_trba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_TBAI[12] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[23]  ( .Q(\pk_scdl_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_bufx1 \REGF/pbmemff41/U1229  ( .Z(\REGF/pbmemff41/n7087 ), .A(
        \REGF/pbmemff41/n7102 ) );
    snl_or02x1 \REGF/pbmemff41/U1246  ( .Z(
        \REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), .A(ph_sa2lt_h), .B(
        \pk_rwrit_h[51] ) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[8]  ( .Q(\pk_sra1_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[8] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[4]  ( .Q(\pk_psae_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[8]  ( .Q(\pk_s45l_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[8]  ( .Q(\pk_sabl_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[1]  ( .Q(\pk_s67l_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[9]  ( .Q(\pk_s89l_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_or02x1 \REGF/pbmemff41/U1247  ( .Z(
        \REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), .A(ph_sa1lt_h), .B(
        \pk_rwrit_h[52] ) );
    snl_and02x1 \REGF/pbmemff41/U1254  ( .Z(\REGF/pbmemff41/RO_PSAS9B551[0] ), 
        .A(ph_lmterr_h), .B(\REGF/pbmemff41/n7103 ) );
    snl_mux21x1 \REGF/pbmemff41/U1261  ( .Z(
        \REGF/pbmemff41/*cell*5493/U75/Z_0 ), .A(PDLIN[19]), .B(\pgldi[3] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[15]  ( .Q(CDOUT[15]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOL[15] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[0]  ( .Q(\REGF/RO_EST1[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(
        \REGF/pbmemff41/RO_PSAS9B551[0] ), .SE(\REGF/pbmemff41/n_2861 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[22]  ( .Q(\REGF/RO_TRCO[26] ), 
        .D(\REGF/pbmemff41/*cell*5493/U61/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7089 ), .SD(\REGF/pbmemff41/RO_TRCOT[22] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[11]  ( .Q(\pk_stdat[11] ), .D(
        \REGF/pbmemff41/*cell*5493/U2/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7099 ), .SD(\REGF/pbmemff41/RO_TRCOT[11] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[2]  ( .Q(\pk_stdat[2] ), .D(
        \REGF/pbmemff41/*cell*5493/U20/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7089 ), .SD(\REGF/pbmemff41/RO_TRCOT[2] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[19]  ( .Q(\pk_sra2_h[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[19] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[19]  ( .Q(\REGF/RO_SRDA[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[19] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[26]  ( .Q(CDOUT[26]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[26] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1268  ( .Z(
        \REGF/pbmemff41/*cell*5493/U61/Z_0 ), .A(PDLIN[26]), .B(\pgldi[10] ), 
        .S(ph_tbllt_h) );
    snl_mux21x1 \REGF/pbmemff41/U1273  ( .Z(
        \REGF/pbmemff41/*cell*5493/U22/DATA2_0 ), .A(PDLIN[1]), .B(\pgldi[1] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[5]  ( .Q(\pk_sra1_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[5] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[5]  ( .Q(\pk_s45l_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[5]  ( .Q(\pk_sabl_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[4]  ( .Q(\pk_s89l_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[22]  ( .Q(CDOUT[22]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOL[22] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[18]  ( .Q(CDOUT[18]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOL[18] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[2]  ( .Q(CDOUT[2]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOL[2] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[23]  ( .Q(\pk_sra1_h[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[23] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[10]  ( .Q(\pk_sra1_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[10] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[27]  ( .Q(\pk_sra2_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_SRA12M[27] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[1]  ( .Q(\pk_scdl_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[14]  ( .Q(\pk_sra2_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[14] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[27]  ( .Q(\REGF/RO_SRDA[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRDA[27] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[14]  ( .Q(\REGF/RO_SRDA[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRDA[14] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOL_reg[11]  ( .Q(CDOUT[11]), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOL[11] ), .SE(
        \pk_rwrit_h[53] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[8]  ( .Q(\pk_scdl_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAE16B_reg[0]  ( .Q(\pk_psae_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[49] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[5]  ( .Q(\pk_s67l_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PSAS9B_reg[4]  ( .Q(\REGF/RO_EST1[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(
        \REGF/pbmemff41/RO_PSAS9B551[4] ), .SE(\REGF/pbmemff41/n_2859 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[15]  ( .Q(\pk_stdat[15] ), .D(
        \REGF/pbmemff41/*cell*5493/U75/Z_0 ), .EN(\REGF/pbmemff41/n8034 ), 
        .RN(\REGF/pbmemff41/n7090 ), .SD(\REGF/pbmemff41/RO_TRCOT[15] ), .SE(
        ph_tblcdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRCOB_reg[6]  ( .Q(\pk_stdat[6] ), .D(
        \REGF/pbmemff41/*cell*5493/U12/DATA2_0 ), .EN(\REGF/pbmemff41/n8035 ), 
        .RN(\REGF/pbmemff41/n7098 ), .SD(\REGF/pbmemff41/RO_TRCOT[6] ), .SE(
        ph_trscdech), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[19]  ( .Q(CDOUT[51]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOH[19] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA128B_reg[19]  ( .Q(\pk_sra1_h[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(
        \REGF/RI_SRA12M[19] ), .SE(\REGF/pbmemff41/*cell*5493/U129/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[4]  ( .Q(\REGF/RO_ERRA[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\pgsadrh[4] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[16]  ( .Q(\pk_trba_h[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(
        \REGF/RI_TBAI[16] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[14]  ( .Q(\pk_scdl_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[5]  ( .Q(\pk_trba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_TBAI[5] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SCDL_reg[27]  ( .Q(\pk_scdl_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[37] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[24]  ( .Q(\pk_s45l_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1260  ( .Z(
        \REGF/pbmemff41/*cell*5493/U77/Z_0 ), .A(PDLIN[18]), .B(\pgldi[2] ), 
        .S(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[19]  ( .Q(\pk_s01l_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[17]  ( .Q(\pk_s45l_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[22]  ( .Q(\pk_sabl_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[11]  ( .Q(\pk_sabl_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[5]  ( .Q(\pk_s01l_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[18]  ( .Q(\pk_s23l_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[25]  ( .Q(\pk_s67l_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[5]  ( .Q(\pk_sefl_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1232  ( .ZN(\REGF/pbmemff41/n7089 ), .A(
        \REGF/pbmemff41/n7087 ) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[2]  ( .Q(\pk_sra2_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[2] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[23]  ( .Q(\REGF/RO_ERRA[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[23] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[16]  ( .Q(\pk_s67l_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[13]  ( .Q(\pk_s89l_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[10]  ( .Q(\REGF/RO_ERRA[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[10] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[20]  ( .Q(\pk_s89l_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[22]  ( .Q(\pk_s23l_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[11]  ( .Q(\pk_s23l_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_and02x1 \REGF/pbmemff41/U1252  ( .Z(\REGF/pbmemff41/RO_PSAS9B551[3] ), 
        .A(ph_lbe2_h), .B(\REGF/pbmemff41/n7103 ) );
    snl_invx05 \REGF/pbmemff41/U1255  ( .ZN(\REGF/pbmemff41/n8037 ), .A(
        ph_trsc_h) );
    snl_mux21x1 \REGF/pbmemff41/U1269  ( .Z(
        \REGF/pbmemff41/*cell*5493/U6/DATA2_0 ), .A(PDLIN[9]), .B(\pgldi[9] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[23]  ( .Q(CDOUT[55]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[23] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[6]  ( .Q(CDOUT[38]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\REGF/RI_PCOH[6] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[19]  ( .Q(\REGF/RO_ERRA[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\pgsadrh[19] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[30]  ( .Q(\pk_s89l_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[29]  ( .Q(\pk_s89l_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[10]  ( .Q(CDOUT[42]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(\REGF/RI_PCOH[10] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[6]  ( .Q(\REGF/RO_SRDA[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_SRDA[6] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[27]  ( .Q(\REGF/RO_ERRA[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[27] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[23]  ( .Q(\pk_s01l_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[10]  ( .Q(\pk_s01l_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[18]  ( .Q(\pk_sabl_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[5]  ( .Q(\pk_s23l_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[25]  ( .Q(\pk_sefl_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[16]  ( .Q(\pk_sefl_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[14]  ( .Q(\REGF/RO_ERRA[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\pgsadrh[14] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[17]  ( .Q(\pk_s89l_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[24]  ( .Q(\pk_s89l_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[27]  ( .Q(CDOUT[59]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOH[27] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[2]  ( .Q(\REGF/RO_SRDA[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[2] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[8]  ( .Q(\pk_trba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(
        \REGF/RI_TBAI[8] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[1]  ( .Q(\pk_trba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(
        \REGF/RI_TBAI[1] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[1]  ( .Q(\pk_s01l_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[1]  ( .Q(\pk_sefl_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[8]  ( .Q(\pk_s23l_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[21]  ( .Q(\pk_s67l_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[12]  ( .Q(\pk_s67l_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[26]  ( .Q(\pk_sabl_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[20]  ( .Q(\pk_s45l_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[15]  ( .Q(\pk_sabl_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[13]  ( .Q(\pk_s45l_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[31]  ( .Q(\pk_sefl_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[28]  ( .Q(\pk_sefl_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[27]  ( .Q(\pk_s01l_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[14]  ( .Q(\pk_s01l_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[30]  ( .Q(\pk_s45l_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[12]  ( .Q(\pk_sefl_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[29]  ( .Q(\pk_s45l_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[21]  ( .Q(\pk_sefl_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[1]  ( .Q(\pk_s23l_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[14]  ( .Q(CDOUT[46]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOH[14] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1272  ( .Z(
        \REGF/pbmemff41/*cell*5493/U24/DATA2_0 ), .A(PDLIN[0]), .B(\pgldi[0] ), 
        .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[2]  ( .Q(CDOUT[34]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[2] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_mux21x1 \REGF/pbmemff41/U1275  ( .Z(
        \REGF/pbmemff41/*cell*5493/U2/DATA2_0 ), .A(PDLIN[11]), .B(\pgldi[11] 
        ), .S(ph_trslt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[6]  ( .Q(\pk_sra2_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRA12M[6] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[15]  ( .Q(\pk_s23l_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[8]  ( .Q(\pk_s01l_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[26]  ( .Q(\pk_s23l_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[8]  ( .Q(\pk_sefl_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[31]  ( .Q(\pk_s67l_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[28]  ( .Q(\pk_s67l_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[25]  ( .Q(CDOUT[57]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7096 ), .SD(\REGF/RI_PCOH[25] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[0]  ( .Q(CDOUT[32]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOH[0] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[4]  ( .Q(\pk_sra2_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[4] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[25]  ( .Q(\pk_s01l_h[25] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[16]  ( .Q(\pk_s01l_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[24]  ( .Q(\pk_s23l_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[17]  ( .Q(\pk_s23l_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[18]  ( .Q(\pk_s45l_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[19]  ( .Q(\pk_s67l_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[23]  ( .Q(\pk_sefl_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[10]  ( .Q(\pk_sefl_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[3]  ( .Q(\pk_s23l_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[16]  ( .Q(CDOUT[48]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOH[16] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[0]  ( .Q(pk_rgbit_h), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_SRDA[0] ), .SE(
        \pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[22]  ( .Q(\pk_s45l_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[24]  ( .Q(\pk_sabl_h[24] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[17]  ( .Q(\pk_sabl_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1235  ( .ZN(\REGF/pbmemff41/n7093 ), .A(
        \REGF/pbmemff41/n7092 ) );
    snl_nand13x1 \REGF/pbmemff41/U1249  ( .ZN(\REGF/pbmemff41/n_2861 ), .A(
        ph_stregwt_h), .B(\REGF/pbmemff41/n8037 ), .C(\REGF/pbmemff41/n7103 )
         );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[9]  ( .Q(CDOUT[41]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(\REGF/RI_PCOH[9] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[9]  ( .Q(\REGF/RO_SRDA[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(
        \REGF/RI_SRDA[9] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[11]  ( .Q(\pk_s45l_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[19]  ( .Q(\pk_sefl_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[3]  ( .Q(\pk_trba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_TBAI[3] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[25]  ( .Q(\REGF/RO_ERRA[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[25] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[15]  ( .Q(\pk_s89l_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[16]  ( .Q(\REGF/RO_ERRA[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[16] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[26]  ( .Q(\pk_s89l_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[3]  ( .Q(\pk_s01l_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[23]  ( .Q(\pk_s67l_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[3]  ( .Q(\pk_sefl_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[21]  ( .Q(CDOUT[53]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\REGF/RI_PCOH[21] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRDA_reg[4]  ( .Q(\REGF/RO_SRDA[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(
        \REGF/RI_SRDA[4] ), .SE(\pk_rwrit_h[50] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[10]  ( .Q(\pk_s67l_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[12]  ( .Q(CDOUT[44]), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(\REGF/RI_PCOH[12] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_PCOH28B_reg[4]  ( .Q(CDOUT[36]), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(\REGF/RI_PCOH[4] ), 
        .SE(\pk_rwrit_h[54] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[0]  ( .Q(\pk_sra2_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_SRA12M[0] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[21]  ( .Q(\pk_s01l_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[12]  ( .Q(\pk_s01l_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[7]  ( .Q(\pk_s23l_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[30]  ( .Q(\pk_sabl_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[29]  ( .Q(\pk_sabl_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[13]  ( .Q(\pk_s23l_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[27]  ( .Q(\pk_sefl_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7098 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[14]  ( .Q(\pk_sefl_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7089 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[20]  ( .Q(\pk_s23l_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff41/U1240  ( .ZN(\REGF/pbmemff41/n7098 ), .A(
        \REGF/pbmemff41/n7097 ) );
    snl_mux21x1 \REGF/pbmemff41/U1267  ( .Z(
        \REGF/pbmemff41/*cell*5493/U63/Z_0 ), .A(PDLIN[25]), .B(\pgldi[9] ), 
        .S(ph_tbllt_h) );
    snl_nor02x1 \REGF/pbmemff41/U1282  ( .ZN(\REGF/pbmemff41/n8034 ), .A(
        \pk_rwrit_h[45] ), .B(ph_tbllt_h) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SRA228B_reg[9]  ( .Q(\pk_sra2_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7093 ), .SD(
        \REGF/RI_SRA12M[9] ), .SE(\REGF/pbmemff41/*cell*5493/U29/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[30]  ( .Q(\pk_s23l_h[30] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7083 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S23L_reg[29]  ( .Q(\pk_s23l_h[29] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[42] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[18]  ( .Q(\pk_s89l_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7090 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[21]  ( .Q(\REGF/RO_ERRA[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7095 ), .SD(\pgsadrh[21] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[7]  ( .Q(\pk_s01l_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SEFL_reg[7]  ( .Q(\pk_sefl_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[36] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[27]  ( .Q(\pk_s67l_h[27] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7101 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S67L_reg[14]  ( .Q(\pk_s67l_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[40] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RRO_ERRA_reg[12]  ( .Q(\REGF/RO_ERRA[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7094 ), .SD(\pgsadrh[12] ), 
        .SE(\pk_rwrit_h[47] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[11]  ( .Q(\pk_s89l_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S89L_reg[22]  ( .Q(\pk_s89l_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7088 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[39] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_TRBA24B_reg[7]  ( .Q(\pk_trba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7085 ), .SD(
        \REGF/RI_TBAI[7] ), .SE(\REGF/pbmemff41/*cell*5493/U27/CONTROL1 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[31]  ( .Q(\pk_s01l_h[31] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7084 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S01L_reg[28]  ( .Q(\pk_s01l_h[28] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7086 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[43] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[26]  ( .Q(\pk_s45l_h[26] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_S45L_reg[15]  ( .Q(\pk_s45l_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7100 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[41] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[20]  ( .Q(\pk_sabl_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7091 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff41/RO_SABL_reg[13]  ( .Q(\pk_sabl_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff41/n7099 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[38] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[16]  ( .Q(\pk_pcs1_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[8]  ( .Q(\pk_pcs1_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[6]  ( .Q(\pk_idcz_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[23]  ( .Q(\pk_saco_lh[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[10]  ( .Q(\pk_saco_lh[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[1]  ( .Q(\pk_pcs1_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[12]  ( .Q(\pk_pcs2_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[20]  ( .Q(\pk_idcx_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[13]  ( .Q(\pk_idcx_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[19]  ( .Q(\pk_saco_lh[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[30]  ( .Q(\REGF/pk_idcx_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[5]  ( .Q(\REGF/pk_scti_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[29]  ( .Q(\REGF/pk_idcx_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[17]  ( .Q(\pk_idcx_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff61/U726  ( .ZN(\REGF/pbmemff61/n6500 ), .A(
        \REGF/pbmemff61/n6502 ) );
    snl_bufx1 \REGF/pbmemff61/U730  ( .Z(\REGF/pbmemff61/n6501 ), .A(
        \REGF/n8052 ) );
    snl_and02x1 \REGF/pbmemff61/U737  ( .Z(\REGF/pbmemff61/RO_EXCO16B882[0] ), 
        .A(\pgbitnoh[0] ), .B(ph_sdirlth) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[12]  ( .Q(\pk_pcs1_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[24]  ( .Q(\REGF/pk_idcx_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[2]  ( .Q(\pk_idcz_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[27]  ( .Q(\pk_saco_hh[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[14]  ( .Q(\pk_saco_lh[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqensnx2 \REGF/pbmemff61/RO_SATI3B_reg[0]  ( .Q(\pk_sati_h[0] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[3] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[5]  ( .Q(\pk_pcs1_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[1]  ( .Q(\REGF/pk_scti_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[16]  ( .Q(\pk_pcs2_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_ERFA1B_reg  ( .Q(\REGF/RO_ERFA[0] ), .D(
        pgperrh), .EN(\REGF/pbmemff61/n6933 ), .RN(\REGF/pbmemff61/n6505 ), 
        .SD(1'b0), .SE(\pk_rwrit_h[0] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[7]  ( .Q(\pk_pcs1_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[3]  ( .Q(\REGF/pk_scti_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[14]  ( .Q(\pk_pcs2_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[9]  ( .Q(\pk_idcz_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_invx1 \REGF/pbmemff61/U731  ( .ZN(\REGF/pbmemff61/n6502 ), .A(
        \REGF/pbmemff61/n6501 ) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[14]  ( .Q(\pk_pcs1_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[10]  ( .Q(\pk_pcs1_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[26]  ( .Q(\REGF/pk_idcx_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[15]  ( .Q(\pk_idcx_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[0]  ( .Q(\pk_idcz_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[25]  ( .Q(\pk_saco_hh[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[16]  ( .Q(\pk_saco_lh[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCSE2B_reg[0]  ( .Q(pk_pcser_h), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[5] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SATI3B_reg[2]  ( .Q(\pk_sati_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[3] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[3]  ( .Q(\pk_pcs1_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[10]  ( .Q(\pk_pcs2_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[7]  ( .Q(\REGF/pk_scti_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[22]  ( .Q(\pk_idcw_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[18]  ( .Q(\pk_idcw_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[22]  ( .Q(\pk_idcx_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[18]  ( .Q(\pk_idcx_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[11]  ( .Q(\pk_idcx_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[4]  ( .Q(\pk_idcz_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[21]  ( .Q(\pk_saco_lh[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[12]  ( .Q(\pk_saco_lh[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_EXCO16B_reg[2]  ( .Q(\REGF/pk_exco_h[2] 
        ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(
        \REGF/pbmemff61/RO_EXCO16B882[2] ), .SE(\REGF/pbmemff61/n_4044 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[11]  ( .Q(\pk_idcw_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[2]  ( .Q(\pk_idcw_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[9]  ( .Q(\pk_idcx_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[20]  ( .Q(\pk_idcz_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[2]  ( .Q(\pk_saco_lh[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[31]  ( .Q(\REGF/pk_idcy_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[28]  ( .Q(\REGF/pk_idcy_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[21]  ( .Q(\pk_idcy_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[13]  ( .Q(\pk_idcz_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[12]  ( .Q(\pk_idcy_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_ARE21B_reg  ( .Q(\REGF/RO_EST2[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[14] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[7]  ( .Q(\pk_idcy_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_and02x1 \REGF/pbmemff61/U736  ( .Z(\REGF/pbmemff61/RO_EXCO16B882[1] ), 
        .A(\pgbitnoh[1] ), .B(ph_sdirlth) );
    snl_or02x1 \REGF/pbmemff61/U738  ( .Z(\REGF/pbmemff61/n_4044 ), .A(
        \pk_rwrit_h[1] ), .B(ph_sdirlth) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[9]  ( .Q(\pk_pcs2_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[4]  ( .Q(\pk_pcs2_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[0]  ( .Q(\pk_idcx_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[25]  ( .Q(\REGF/pk_idcy_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[30]  ( .Q(\REGF/pk_idcz_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[29]  ( .Q(\REGF/pk_idcz_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SRE21B_reg  ( .Q(\REGF/RO_EST2[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[16] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[16]  ( .Q(\pk_idcy_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[24]  ( .Q(\REGF/pk_idcz_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[6]  ( .Q(\pk_saco_lh[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[17]  ( .Q(\pk_idcz_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[0]  ( .Q(\pk_pcs2_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[26]  ( .Q(\REGF/pk_idcw_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[15]  ( .Q(\pk_idcw_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[4]  ( .Q(\pk_idcx_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SASE4B_reg[3]  ( .Q(pk_sasea_h), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[4] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[6]  ( .Q(\pk_idcw_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[3]  ( .Q(\pk_idcy_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[2]  ( .Q(\pk_pcs2_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[4]  ( .Q(\pk_idcw_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[1]  ( .Q(\pk_idcy_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_ARE31B_reg  ( .Q(\REGF/RO_EST2[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[13] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[6]  ( .Q(\pk_idcx_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[24]  ( .Q(\REGF/pk_idcw_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[17]  ( .Q(\pk_idcw_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SASE4B_reg[1]  ( .Q(\pk_saseo_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[4] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[20]  ( .Q(\pk_idcw_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[13]  ( .Q(\pk_idcw_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[27]  ( .Q(\REGF/pk_idcy_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[8]  ( .Q(\pk_idcy_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[26]  ( .Q(\REGF/pk_idcz_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[15]  ( .Q(\pk_idcz_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[4]  ( .Q(\pk_saco_lh[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[14]  ( .Q(\pk_idcy_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[6]  ( .Q(\pk_pcs2_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[18]  ( .Q(\pk_idcz_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[30]  ( .Q(\REGF/pk_idcw_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[9]  ( .Q(\pk_idcw_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[0]  ( .Q(\pk_idcw_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[2]  ( .Q(\pk_idcx_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[19]  ( .Q(\pk_idcy_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[9]  ( .Q(\pk_saco_lh[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[23]  ( .Q(\pk_idcy_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[5]  ( .Q(\pk_idcy_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[10]  ( .Q(\pk_idcy_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_EXCO16B_reg[0]  ( .Q(\REGF/pk_exco_h[0] 
        ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(
        \REGF/pbmemff61/RO_EXCO16B882[0] ), .SE(\REGF/pbmemff61/n_4044 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[29]  ( .Q(\REGF/pk_idcw_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[7]  ( .Q(\pk_pcs2_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[21]  ( .Q(\pk_idcw_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[12]  ( .Q(\pk_idcw_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[22]  ( .Q(\pk_idcz_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[0]  ( .Q(\pk_saco_lh[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[11]  ( .Q(\pk_idcz_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[3]  ( .Q(\pk_idcx_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[19]  ( .Q(\pk_idcz_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff61/U727  ( .ZN(\REGF/pbmemff61/n6506 ), .A(
        \REGF/pbmemff61/n6502 ) );
    snl_invx2 \REGF/pbmemff61/U728  ( .ZN(\REGF/pbmemff61/n6504 ), .A(
        \REGF/pbmemff61/n6502 ) );
    snl_invx05 \REGF/pbmemff61/U733  ( .ZN(\REGF/pbmemff61/n6933 ), .A(
        ph_cperlt_h) );
    snl_and02x1 \REGF/pbmemff61/U734  ( .Z(\REGF/pbmemff61/RO_EXCO16B882[3] ), 
        .A(\pgbitnoh[3] ), .B(ph_sdirlth) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[3]  ( .Q(\pk_pcs2_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[31]  ( .Q(\REGF/pk_idcw_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[28]  ( .Q(\REGF/pk_idcw_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[8]  ( .Q(\pk_idcw_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[1]  ( .Q(\pk_idcw_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[18]  ( .Q(\pk_idcy_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[8]  ( .Q(\pk_saco_lh[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[4]  ( .Q(\pk_idcy_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[22]  ( .Q(\pk_idcy_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[11]  ( .Q(\pk_idcy_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[5]  ( .Q(\pk_idcw_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[23]  ( .Q(\pk_idcz_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[1]  ( .Q(\pk_saco_lh[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_EXCO16B_reg[1]  ( .Q(\REGF/pk_exco_h[1] 
        ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(
        \REGF/pbmemff61/RO_EXCO16B882[1] ), .SE(\REGF/pbmemff61/n_4044 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[10]  ( .Q(\pk_idcz_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[0]  ( .Q(\pk_idcy_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SASE4B_reg[0]  ( .Q(pk_sased_h), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[4] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[25]  ( .Q(\REGF/pk_idcw_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[16]  ( .Q(\pk_idcw_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[7]  ( .Q(\pk_idcx_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[27]  ( .Q(\REGF/pk_idcz_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[14]  ( .Q(\pk_idcz_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[5]  ( .Q(\pk_saco_lh[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[26]  ( .Q(\REGF/pk_idcy_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[9]  ( .Q(\pk_idcy_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[15]  ( .Q(\pk_idcy_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[8]  ( .Q(\pk_pcs2_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[24]  ( .Q(\REGF/pk_idcy_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[17]  ( .Q(\pk_idcy_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[25]  ( .Q(\REGF/pk_idcz_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[7]  ( .Q(\pk_saco_lh[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[16]  ( .Q(\pk_idcz_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[1]  ( .Q(\pk_pcs2_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[5]  ( .Q(\pk_idcx_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SASE4B_reg[2]  ( .Q(\pk_saseo_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[4] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[27]  ( .Q(\REGF/pk_idcw_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[14]  ( .Q(\pk_idcw_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[7]  ( .Q(\pk_idcw_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[2]  ( .Q(\pk_idcy_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_STIM1B_reg  ( .Q(\REGF/RO_PSTA[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[18] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff61/U729  ( .ZN(\REGF/pbmemff61/n6505 ), .A(
        \REGF/pbmemff61/n6502 ) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[15]  ( .Q(\pk_pcs1_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[5]  ( .Q(\pk_pcs2_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[23]  ( .Q(\pk_idcw_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[19]  ( .Q(\pk_idcw_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_EXCO16B_reg[3]  ( .Q(\REGF/pk_exco_h[3] 
        ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(
        \REGF/pbmemff61/RO_EXCO16B882[3] ), .SE(\REGF/pbmemff61/n_4044 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[10]  ( .Q(\pk_idcw_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCW_reg[3]  ( .Q(\pk_idcw_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[10] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[8]  ( .Q(\pk_idcx_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[21]  ( .Q(\pk_idcz_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[3]  ( .Q(\pk_saco_lh[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[30]  ( .Q(\REGF/pk_idcy_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[20]  ( .Q(\pk_idcy_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[12]  ( .Q(\pk_idcz_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[13]  ( .Q(\pk_idcy_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[29]  ( .Q(\REGF/pk_idcy_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCY_reg[6]  ( .Q(\pk_idcy_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[8] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[1]  ( .Q(\pk_idcx_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[31]  ( .Q(\REGF/pk_idcz_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[28]  ( .Q(\REGF/pk_idcz_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCSE2B_reg[1]  ( .Q(pk_pcsee_h), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[5] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff61/U732  ( .ZN(\REGF/pbmemff61/n6503 ), .A(
        \REGF/pbmemff61/n6502 ) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[2]  ( .Q(\pk_pcs1_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[19]  ( .Q(\pk_idcx_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[6]  ( .Q(\REGF/pk_scti_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[18]  ( .Q(\pk_pcs2_h[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[11]  ( .Q(\pk_pcs2_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[5]  ( .Q(\pk_idcz_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[20]  ( .Q(\pk_saco_lh[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[13]  ( .Q(\pk_saco_lh[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[23]  ( .Q(\pk_idcx_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[10]  ( .Q(\pk_idcx_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[18]  ( .Q(\pk_pcs1_h[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[11]  ( .Q(\pk_pcs1_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[6]  ( .Q(\pk_pcs1_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[15]  ( .Q(\pk_pcs2_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[2]  ( .Q(\REGF/pk_scti_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[8]  ( .Q(\pk_idcz_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SRAS1B_reg  ( .Q(\REGF/RO_EST2[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[19] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[13]  ( .Q(\pk_pcs1_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[27]  ( .Q(\REGF/pk_idcx_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[14]  ( .Q(\pk_idcx_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[25]  ( .Q(\REGF/pk_idcx_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[16]  ( .Q(\pk_idcx_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[1]  ( .Q(\pk_idcz_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[24]  ( .Q(\pk_saco_hh[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[17]  ( .Q(\pk_saco_lh[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[3]  ( .Q(\pk_idcz_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqensnx2 \REGF/pbmemff61/RO_SATI3B_reg[1]  ( .Q(\pk_sati_h[1] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[3] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[26]  ( .Q(\pk_saco_hh[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[15]  ( .Q(\pk_saco_lh[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_ARE11B_reg  ( .Q(\REGF/RO_EST2[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[15] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[4]  ( .Q(\pk_pcs1_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[17]  ( .Q(\pk_pcs2_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[0]  ( .Q(\REGF/pk_scti_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_and02x1 \REGF/pbmemff61/U735  ( .Z(\REGF/pbmemff61/RO_EXCO16B882[2] ), 
        .A(\pgbitnoh[2] ), .B(ph_sdirlth) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[17]  ( .Q(\pk_pcs1_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[9]  ( .Q(\pk_pcs1_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6503 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[12]  ( .Q(\pk_idcx_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCZ_reg[7]  ( .Q(\pk_idcz_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[7] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[22]  ( .Q(\pk_saco_lh[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[11]  ( .Q(\pk_saco_lh[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SRE11B_reg  ( .Q(\REGF/RO_PSTA[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[17] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS119B_reg[0]  ( .Q(\pk_pcs1_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[12] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[31]  ( .Q(\REGF/pk_idcx_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6505 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[28]  ( .Q(\REGF/pk_idcx_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6504 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_IDCX_reg[21]  ( .Q(\pk_idcx_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6501 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[9] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SACO28B_reg[18]  ( .Q(\pk_saco_lh[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6506 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[6] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_SCTI8B_reg[4]  ( .Q(\REGF/pk_scti_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[2] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff61/RO_PCS219B_reg[13]  ( .Q(\pk_pcs2_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff61/n6500 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[11] ), .CP(SCLK) );
    snl_aoi223x0 \CONS/gte_124/U6  ( .ZN(\CONS/gte_124/n15 ), .A(
        \CONS/gte_124/n16 ), .B(\CONS/gte_124/n17 ), .C(\CONS/gte_124/n18 ), 
        .D(\pk_pc_h[16] ), .E(\CONS/gte_124/n19 ), .F(\pk_pc_h[17] ), .G(
        \CONS/gte_124/n24 ) );
    snl_nor02x1 \CONS/gte_124/U14  ( .ZN(\CONS/gte_124/n47 ), .A(\pk_pc_h[9] ), 
        .B(\CONS/gte_124/n43 ) );
    snl_invx05 \CONS/gte_124/U21  ( .ZN(\CONS/gte_124/n29 ), .A(\pk_pcs1_h[1] 
        ) );
    snl_invx05 \CONS/gte_124/U28  ( .ZN(\CONS/gte_124/n43 ), .A(\pk_pcs1_h[9] 
        ) );
    snl_invx05 \CONS/gte_124/U33  ( .ZN(\CONS/gte_124/n55 ), .A(\pk_pc_h[14] )
         );
    snl_oai023x0 \CONS/gte_124/U7  ( .ZN(\CONS/n298 ), .A(\CONS/gte_124/n25 ), 
        .B(\CONS/gte_124/n15 ), .C(\CONS/gte_124/n26 ), .D(\pk_pcs1_h[18] ), 
        .E(\CONS/gte_124/n27 ) );
    snl_aoi1b12x0 \CONS/gte_124/U8  ( .ZN(\CONS/gte_124/n28 ), .A(\pk_pc_h[1] 
        ), .B(\CONS/gte_124/n29 ), .C(\pk_pcs1_h[0] ), .D(\pk_pc_h[0] ) );
    snl_and02x1 \CONS/gte_124/U13  ( .Z(\CONS/gte_124/n45 ), .A(
        \CONS/gte_124/n46 ), .B(\pk_pcs1_h[10] ) );
    snl_invx05 \CONS/gte_124/U34  ( .ZN(\CONS/gte_124/n61 ), .A(\pk_pc_h[15] )
         );
    snl_nand02x1 \CONS/gte_124/U41  ( .ZN(\CONS/gte_124/n33 ), .A(
        \pk_pcs1_h[3] ), .B(\CONS/gte_124/n58 ) );
    snl_nand12x1 \CONS/gte_124/U46  ( .ZN(\CONS/gte_124/n49 ), .A(
        \pk_pc_h[12] ), .B(\pk_pcs1_h[12] ) );
    snl_invx05 \CONS/gte_124/U26  ( .ZN(\CONS/gte_124/n59 ), .A(\pk_pc_h[7] )
         );
    snl_oai223x0 \CONS/gte_124/U48  ( .ZN(\CONS/gte_124/n17 ), .A(
        \CONS/gte_124/n56 ), .B(\CONS/gte_124/n48 ), .C(\CONS/gte_124/n54 ), 
        .D(\pk_pcs1_h[14] ), .E(\CONS/gte_124/n55 ), .F(\pk_pcs1_h[15] ), .G(
        \CONS/gte_124/n61 ) );
    snl_aoi223x0 \CONS/gte_124/U9  ( .ZN(\CONS/gte_124/n30 ), .A(
        \CONS/gte_124/n31 ), .B(\CONS/gte_124/n32 ), .C(\CONS/gte_124/n33 ), 
        .D(\pk_pc_h[5] ), .E(\CONS/gte_124/n34 ), .F(\pk_pc_h[4] ), .G(
        \CONS/gte_124/n35 ) );
    snl_aoi223x0 \CONS/gte_124/U12  ( .ZN(\CONS/gte_124/n39 ), .A(
        \CONS/gte_124/n40 ), .B(\CONS/gte_124/n41 ), .C(\CONS/gte_124/n42 ), 
        .D(\pk_pc_h[9] ), .E(\CONS/gte_124/n43 ), .F(\pk_pc_h[8] ), .G(
        \CONS/gte_124/n44 ) );
    snl_invx05 \CONS/gte_124/U35  ( .ZN(\CONS/gte_124/n19 ), .A(
        \pk_pcs1_h[16] ) );
    snl_invx05 \CONS/gte_124/U27  ( .ZN(\CONS/gte_124/n44 ), .A(\pk_pcs1_h[8] 
        ) );
    snl_nand12x1 \CONS/gte_124/U40  ( .ZN(\CONS/gte_124/n31 ), .A(\pk_pc_h[4] 
        ), .B(\pk_pcs1_h[4] ) );
    snl_invx05 \CONS/gte_124/U20  ( .ZN(\CONS/gte_124/n57 ), .A(\pk_pcs1_h[2] 
        ) );
    snl_nand12x1 \CONS/gte_124/U49  ( .ZN(\CONS/gte_124/n16 ), .A(
        \pk_pc_h[16] ), .B(\pk_pcs1_h[16] ) );
    snl_invx05 \CONS/gte_124/U29  ( .ZN(\CONS/gte_124/n46 ), .A(\pk_pc_h[10] )
         );
    snl_nand02x1 \CONS/gte_124/U47  ( .ZN(\CONS/gte_124/n51 ), .A(
        \pk_pcs1_h[11] ), .B(\CONS/gte_124/n60 ) );
    snl_and02x1 \CONS/gte_124/U10  ( .Z(\CONS/gte_124/n36 ), .A(
        \CONS/gte_124/n37 ), .B(\pk_pcs1_h[6] ) );
    snl_aoi223x0 \CONS/gte_124/U15  ( .ZN(\CONS/gte_124/n48 ), .A(
        \CONS/gte_124/n49 ), .B(\CONS/gte_124/n50 ), .C(\CONS/gte_124/n51 ), 
        .D(\pk_pc_h[13] ), .E(\CONS/gte_124/n52 ), .F(\pk_pc_h[12] ), .G(
        \CONS/gte_124/n53 ) );
    snl_nor02x1 \CONS/gte_124/U17  ( .ZN(\CONS/gte_124/n56 ), .A(\pk_pc_h[13] 
        ), .B(\CONS/gte_124/n52 ) );
    snl_invx05 \CONS/gte_124/U22  ( .ZN(\CONS/gte_124/n58 ), .A(\pk_pc_h[3] )
         );
    snl_invx05 \CONS/gte_124/U32  ( .ZN(\CONS/gte_124/n52 ), .A(
        \pk_pcs1_h[13] ) );
    snl_ao2b2b2x0 \CONS/gte_124/U39  ( .Z(\CONS/gte_124/n32 ), .A(
        \pk_pcs1_h[3] ), .B(\CONS/gte_124/n58 ), .C(\CONS/gte_124/n28 ), .D(
        \CONS/gte_124/n62 ), .E(\CONS/gte_124/n57 ), .F(\pk_pc_h[2] ) );
    snl_invx05 \CONS/gte_124/U30  ( .ZN(\CONS/gte_124/n60 ), .A(\pk_pc_h[11] )
         );
    snl_oai223x0 \CONS/gte_124/U42  ( .ZN(\CONS/gte_124/n41 ), .A(
        \CONS/gte_124/n38 ), .B(\CONS/gte_124/n30 ), .C(\CONS/gte_124/n36 ), 
        .D(\pk_pcs1_h[6] ), .E(\CONS/gte_124/n37 ), .F(\pk_pcs1_h[7] ), .G(
        \CONS/gte_124/n59 ) );
    snl_oai223x0 \CONS/gte_124/U45  ( .ZN(\CONS/gte_124/n50 ), .A(
        \CONS/gte_124/n47 ), .B(\CONS/gte_124/n39 ), .C(\CONS/gte_124/n45 ), 
        .D(\pk_pcs1_h[10] ), .E(\CONS/gte_124/n46 ), .F(\pk_pcs1_h[11] ), .G(
        \CONS/gte_124/n60 ) );
    snl_nor02x1 \CONS/gte_124/U11  ( .ZN(\CONS/gte_124/n38 ), .A(\pk_pc_h[5] ), 
        .B(\CONS/gte_124/n34 ) );
    snl_nor02x1 \CONS/gte_124/U19  ( .ZN(\CONS/gte_124/n25 ), .A(\pk_pc_h[17] 
        ), .B(\CONS/gte_124/n24 ) );
    snl_invx05 \CONS/gte_124/U25  ( .ZN(\CONS/gte_124/n37 ), .A(\pk_pc_h[6] )
         );
    snl_invx05 \CONS/gte_124/U37  ( .ZN(\CONS/gte_124/n27 ), .A(\pk_pc_h[18] )
         );
    snl_nand02x1 \CONS/gte_124/U50  ( .ZN(\CONS/gte_124/n18 ), .A(
        \pk_pcs1_h[15] ), .B(\CONS/gte_124/n61 ) );
    snl_and02x1 \CONS/gte_124/U16  ( .Z(\CONS/gte_124/n54 ), .A(
        \CONS/gte_124/n55 ), .B(\pk_pcs1_h[14] ) );
    snl_and02x1 \CONS/gte_124/U18  ( .Z(\CONS/gte_124/n26 ), .A(
        \CONS/gte_124/n27 ), .B(\pk_pcs1_h[18] ) );
    snl_invx05 \CONS/gte_124/U36  ( .ZN(\CONS/gte_124/n24 ), .A(
        \pk_pcs1_h[17] ) );
    snl_nand12x1 \CONS/gte_124/U43  ( .ZN(\CONS/gte_124/n40 ), .A(\pk_pc_h[8] 
        ), .B(\pk_pcs1_h[8] ) );
    snl_invx05 \CONS/gte_124/U23  ( .ZN(\CONS/gte_124/n35 ), .A(\pk_pcs1_h[4] 
        ) );
    snl_invx05 \CONS/gte_124/U24  ( .ZN(\CONS/gte_124/n34 ), .A(\pk_pcs1_h[5] 
        ) );
    snl_invx05 \CONS/gte_124/U31  ( .ZN(\CONS/gte_124/n53 ), .A(
        \pk_pcs1_h[12] ) );
    snl_oai022x1 \CONS/gte_124/U38  ( .ZN(\CONS/gte_124/n62 ), .A(\pk_pc_h[1] 
        ), .B(\CONS/gte_124/n29 ), .C(\pk_pc_h[2] ), .D(\CONS/gte_124/n57 ) );
    snl_nand02x1 \CONS/gte_124/U44  ( .ZN(\CONS/gte_124/n42 ), .A(
        \pk_pcs1_h[7] ), .B(\CONS/gte_124/n59 ) );
    snl_ao123x1 \CODEIF/CNT/U185  ( .Z(\CODEIF/CNT/wpfcen ), .A(st_cfctl), .B(
        \CODEIF/CNT/n3805 ), .C(\CODEIF/CNT/n3806 ), .D(\CODEIF/CNT/n3768 ), 
        .E(\CODEIF/CNT/n3804 ), .F(\CODEIF/CNT/n3807 ) );
    snl_nand14x0 \CODEIF/CNT/U191  ( .ZN(\CODEIF/CNT/nst[2] ), .A(
        \CODEIF/CNT/n3779 ), .B(\CODEIF/CNT/n3780 ), .C(\CODEIF/CNT/n3781 ), 
        .D(\CODEIF/CNT/n3782 ) );
    snl_aoi013x0 \CODEIF/CNT/U198  ( .ZN(\CODEIF/CNT/n3787 ), .A(st_cfctl), 
        .B(\CODEIF/CNT/n3803 ), .C(\CODEIF/CNT/n3804 ), .D(\CODEIF/CNT/n3771 )
         );
    snl_aoi012x1 \CODEIF/CNT/U204  ( .ZN(\CODEIF/CNT/n3815 ), .A(
        \CODEIF/CNT/n3803 ), .B(\CODEIF/CNT/n3805 ), .C(\CODEIF/CNT/n3816 ) );
    snl_nand02x1 \CODEIF/CNT/U223  ( .ZN(\CODEIF/CNT/n3799 ), .A(
        \CODEIF/write_prtect ), .B(cif_byte) );
    snl_nor02x1 \CODEIF/CNT/U238  ( .ZN(\CODEIF/CNT/n3830 ), .A(
        \CODEIF/CNT/n3836 ), .B(\CODEIF/CNT/n3807 ) );
    snl_invx05 \CODEIF/CNT/U256  ( .ZN(\CODEIF/CNT/n3783 ), .A(
        \CODEIF/CNT/wwbregen ) );
    snl_invx05 \CODEIF/CNT/U271  ( .ZN(\CODEIF/CNT/n3789 ), .A(
        \CODEIF/CNT/n3802 ) );
    snl_nor02x1 \CODEIF/CNT/U196  ( .ZN(\CODEIF/friend_in ), .A(cf_wait), .B(
        \CODEIF/CNT/n3796 ) );
    snl_nand02x1 \CODEIF/CNT/U211  ( .ZN(\CODEIF/CNT/n3794 ), .A(
        \CODEIF/CNT/cst[3] ), .B(\CODEIF/CNT/n3818 ) );
    snl_invx05 \CODEIF/CNT/U216  ( .ZN(\CODEIF/CNT/n3821 ), .A(
        \CODEIF/CNT/cst[1] ) );
    snl_xor2x0 \CODEIF/CNT/U231  ( .Z(\CODEIF/CNT/n3831 ), .A(st_cfctl), .B(
        cif_cont) );
    snl_oai223x0 \CODEIF/CNT/U244  ( .ZN(\CODEIF/CNT/n3775 ), .A(
        \CODEIF/CNT/n3839 ), .B(\CODEIF/fm_config[1] ), .C(
        \CODEIF/fm_config[0] ), .D(\CODEIF/CNT/n3825 ), .E(\CODEIF/CNT/n3776 ), 
        .F(cf_wait), .G(\CODEIF/CNT/n3840 ) );
    snl_invx05 \CODEIF/CNT/U263  ( .ZN(\CODEIF/CNT/n3804 ), .A(
        \CODEIF/CNT/n3822 ) );
    snl_nor02x1 \CODEIF/CNT/U236  ( .ZN(\CODEIF/CNT/n3811 ), .A(cif_byte), .B(
        cif_cont) );
    snl_aoi122x0 \CODEIF/CNT/U243  ( .ZN(\CODEIF/CNT/n3778 ), .A(
        \CODEIF/CNT/n3827 ), .B(\CODEIF/CNT/n3814 ), .C(\CODEIF/CNT/n3833 ), 
        .D(\CODEIF/CNT/n3825 ), .E(\CODEIF/CNT/n3779 ) );
    snl_nor03x0 \CODEIF/CNT/U258  ( .ZN(\CODEIF/wprotect1 ), .A(
        \CODEIF/CNT/n3790 ), .B(\CODEIF/write_prtect ), .C(\CODEIF/CNT/n3820 )
         );
    snl_invx05 \CODEIF/CNT/U264  ( .ZN(\CODEIF/CNT/n3767 ), .A(
        \CODEIF/CNT/n3794 ) );
    snl_oai122x0 \CODEIF/CNT/U197  ( .ZN(\CODEIF/frpend_in ), .A(
        \CODEIF/CNT/n3797 ), .B(\CODEIF/CNT/n3798 ), .C(\CODEIF/CNT/n3790 ), 
        .D(\CODEIF/CNT/n3799 ), .E(\CODEIF/CNT/n3800 ) );
    snl_nand02x1 \CODEIF/CNT/U203  ( .ZN(\CODEIF/CNT/n3814 ), .A(
        \CODEIF/CNT/cst[4] ), .B(\CODEIF/CNT/cst[3] ) );
    snl_nand02x1 \CODEIF/CNT/U218  ( .ZN(\CODEIF/CNT/n3823 ), .A(
        \CODEIF/CNT/cst[0] ), .B(\CODEIF/CNT/cst[2] ) );
    snl_nor02x1 \CODEIF/CNT/U251  ( .ZN(\CODEIF/CNT/n3836 ), .A(
        \CODEIF/CNT/n3797 ), .B(\CODEIF/CNT/n3822 ) );
    snl_nand02x1 \CODEIF/CNT/U276  ( .ZN(\CODEIF/CNT/n3780 ), .A(
        \CODEIF/fm_config[1] ), .B(\CODEIF/CNT/n3841 ) );
    snl_nand03x0 \CODEIF/CNT/U224  ( .ZN(\CODEIF/CNT/n3777 ), .A(
        \CODEIF/CNT/n3804 ), .B(\CODEIF/CNT/n3810 ), .C(\CODEIF/CNT/cst[0] )
         );
    snl_nor02x1 \CODEIF/CNT/U202  ( .ZN(\CODEIF/CNT/n3766 ), .A(
        \CODEIF/CNT/cst[2] ), .B(\CODEIF/CNT/n3809 ) );
    snl_invx05 \CODEIF/CNT/U210  ( .ZN(\CODEIF/CNT/n3820 ), .A(cif_byte) );
    snl_aoi113x0 \CODEIF/CNT/U242  ( .ZN(\CODEIF/CNT/n3782 ), .A(
        \CODEIF/CNT/cst[1] ), .B(\CODEIF/CNT/n3809 ), .C(\CODEIF/CNT/n3838 ), 
        .D(\CODEIF/CNT/n3816 ), .E(\CODEIF/CNT/n3772 ) );
    snl_invx05 \CODEIF/CNT/U265  ( .ZN(\CODEIF/CNT/n3829 ), .A(
        \CODEIF/CNT/n3827 ) );
    snl_nor03x0 \CODEIF/CNT/U259  ( .ZN(\CODEIF/CNT/n3793 ), .A(
        \CODEIF/CNT/n3768 ), .B(st_cfctl), .C(\CODEIF/CNT/n3822 ) );
    snl_ffqrnx1 \CODEIF/CNT/cst_reg[0]  ( .Q(\CODEIF/CNT/cst[0] ), .D(
        \CODEIF/CNT/nst[0] ), .RN(\CODEIF/n3862 ), .CP(SCLK) );
    snl_nand02x1 \CODEIF/CNT/U237  ( .ZN(\CODEIF/CNT/n3828 ), .A(cif_byte), 
        .B(\CODEIF/CNT/n3835 ) );
    snl_nor02x1 \CODEIF/CNT/U225  ( .ZN(\CODEIF/CNT/n3827 ), .A(
        \CODEIF/CNT/n3821 ), .B(\CODEIF/CNT/cst[2] ) );
    snl_ffqrnx1 \CODEIF/CNT/cst_reg[4]  ( .Q(\CODEIF/CNT/cst[4] ), .D(
        \CODEIF/CNT/nst[4] ), .RN(\CODEIF/n3862 ), .CP(SCLK) );
    snl_aoi112x0 \CODEIF/CNT/U250  ( .ZN(\CODEIF/CNT/n3771 ), .A(
        \CODEIF/CNT/n3808 ), .B(\CODEIF/CNT/n3823 ), .C(\CODEIF/CNT/cst[1] ), 
        .D(\CODEIF/CNT/n3822 ) );
    snl_nand03x0 \CODEIF/CNT/U277  ( .ZN(\CODEIF/CNT/n3832 ), .A(
        \CODEIF/CNT/n3819 ), .B(\CODEIF/CNT/n3820 ), .C(cif_cont) );
    snl_oai112x2 \CODEIF/CNT/U186  ( .ZN(\CODEIF/fadren ), .A(
        \CODEIF/CNT/n3801 ), .B(\CODEIF/CNT/n3802 ), .C(\CODEIF/CNT/n3783 ), 
        .D(\CODEIF/CNT/n3786 ) );
    snl_oai012x1 \CODEIF/CNT/U187  ( .ZN(pgrstith), .A(\CODEIF/CNT/cst[1] ), 
        .B(\CODEIF/CNT/n3766 ), .C(\CODEIF/CNT/n3767 ) );
    snl_or08x1 \CODEIF/CNT/U189  ( .Z(\CODEIF/CNT/nst[0] ), .A(
        \CODEIF/CNT/n3769 ), .B(\CODEIF/CNT/n3770 ), .C(\CODEIF/CNT/n3771 ), 
        .D(\CODEIF/CNT/wwbregen ), .E(\CODEIF/CNT/n3772 ), .F(
        \CODEIF/CNT/n3773 ), .G(\CODEIF/CNT/n3774 ), .H(\CODEIF/CNT/n3775 ) );
    snl_nand14x0 \CODEIF/CNT/U190  ( .ZN(\CODEIF/CNT/nst[1] ), .A(
        \CODEIF/CNT/n3769 ), .B(\CODEIF/CNT/n3776 ), .C(\CODEIF/CNT/n3777 ), 
        .D(\CODEIF/CNT/n3778 ) );
    snl_nand12x1 \CODEIF/CNT/U199  ( .ZN(\CODEIF/CNT/n3808 ), .A(
        \CODEIF/CNT/cst[2] ), .B(\CODEIF/CNT/n3809 ) );
    snl_nor02x1 \CODEIF/CNT/U205  ( .ZN(\CODEIF/CNT/n3810 ), .A(
        \CODEIF/CNT/cst[1] ), .B(\CODEIF/CNT/cst[2] ) );
    snl_nor02x1 \CODEIF/CNT/U219  ( .ZN(\CODEIF/CNT/n3824 ), .A(
        \CODEIF/CNT/n3823 ), .B(\CODEIF/CNT/cst[4] ) );
    snl_nand02x1 \CODEIF/CNT/U222  ( .ZN(\CODEIF/CNT/n3798 ), .A(
        \CODEIF/CNT/n3805 ), .B(\CODEIF/CNT/n3818 ) );
    snl_aoi123x0 \CODEIF/CNT/U239  ( .ZN(\CODEIF/CNT/n3788 ), .A(st_cfctl), 
        .B(\CODEIF/CNT/n3819 ), .C(\CODEIF/CNT/n3811 ), .D(\CODEIF/CNT/n3827 ), 
        .E(\CODEIF/CNT/n3804 ), .F(\CODEIF/CNT/n3779 ) );
    snl_nor02x1 \CODEIF/CNT/U257  ( .ZN(\CODEIF/wprotect0 ), .A(
        \CODEIF/CNT/n3768 ), .B(\CODEIF/CNT/n3794 ) );
    snl_invx05 \CODEIF/CNT/U270  ( .ZN(\CODEIF/CNT/n3812 ), .A(
        \CODEIF/CNT/n3797 ) );
    snl_nand03x0 \CODEIF/CNT/U217  ( .ZN(\CODEIF/CNT/n3797 ), .A(
        \CODEIF/CNT/cst[2] ), .B(\CODEIF/CNT/n3809 ), .C(\CODEIF/CNT/cst[1] )
         );
    snl_nand02x1 \CODEIF/CNT/U230  ( .ZN(\CODEIF/CNT/n3802 ), .A(
        \CODEIF/CNT/n3831 ), .B(\CODEIF/CNT/n3820 ) );
    snl_invx05 \CODEIF/CNT/U245  ( .ZN(\CODEIF/CNT/n3790 ), .A(
        \CODEIF/CNT/n3819 ) );
    snl_nor02x1 \CODEIF/CNT/U262  ( .ZN(\CODEIF/CNT/n3813 ), .A(
        \CODEIF/CNT/n3777 ), .B(\CODEIF/CNT/n3825 ) );
    snl_ffqrnx1 \CODEIF/CNT/cst_reg[2]  ( .Q(\CODEIF/CNT/cst[2] ), .D(
        \CODEIF/CNT/nst[2] ), .RN(\CODEIF/n3862 ), .CP(SCLK) );
    snl_nand04x0 \CODEIF/CNT/U192  ( .ZN(\CODEIF/CNT/nst[3] ), .A(
        \CODEIF/CNT/n3783 ), .B(\CODEIF/CNT/n3776 ), .C(\CODEIF/CNT/n3784 ), 
        .D(\CODEIF/CNT/n3785 ) );
    snl_nand02x1 \CODEIF/CNT/U207  ( .ZN(\CODEIF/CNT/n3801 ), .A(
        \CODEIF/CNT/n3817 ), .B(\CODEIF/CNT/n3809 ) );
    snl_nand02x1 \CODEIF/CNT/U220  ( .ZN(\CODEIF/CNT/n3825 ), .A(
        \CODEIF/fm_config[1] ), .B(\CODEIF/fm_config[0] ) );
    snl_nor02x1 \CODEIF/CNT/U255  ( .ZN(\CODEIF/CNT/wwbregen ), .A(
        \CODEIF/CNT/n3805 ), .B(\CODEIF/CNT/n3801 ) );
    snl_invx05 \CODEIF/CNT/U269  ( .ZN(\CODEIF/wpfcinc ), .A(
        \CODEIF/CNT/n3787 ) );
    snl_nor03x0 \CODEIF/CNT/U272  ( .ZN(\CODEIF/CNT/n3840 ), .A(
        \CODEIF/CNT/n3807 ), .B(\CODEIF/CNT/n3836 ), .C(\CODEIF/CNT/n3813 ) );
    snl_ffqrnx1 \CODEIF/CNT/cst_reg[3]  ( .Q(\CODEIF/CNT/cst[3] ), .D(
        \CODEIF/CNT/nst[3] ), .RN(\CODEIF/n3862 ), .CP(SCLK) );
    snl_invx05 \CODEIF/CNT/U215  ( .ZN(\CODEIF/CNT/n3809 ), .A(
        \CODEIF/CNT/cst[0] ) );
    snl_nand03x0 \CODEIF/CNT/U229  ( .ZN(\CODEIF/CNT/n3776 ), .A(
        \CODEIF/CNT/cst[3] ), .B(\CODEIF/CNT/n3817 ), .C(\CODEIF/CNT/cst[0] )
         );
    snl_nor03x0 \CODEIF/CNT/U247  ( .ZN(\CODEIF/CNT/n3770 ), .A(
        \CODEIF/CNT/n3821 ), .B(\CODEIF/CNT/n3805 ), .C(\CODEIF/CNT/n3791 ) );
    snl_nor02x1 \CODEIF/CNT/U260  ( .ZN(\CODEIF/CNT/n3772 ), .A(
        \CODEIF/CNT/n3798 ), .B(\CODEIF/CNT/n3768 ) );
    snl_muxi21x1 \CODEIF/CNT/U232  ( .ZN(\CODEIF/CNT/n3774 ), .A(
        \CODEIF/CNT/n3832 ), .B(\CODEIF/CNT/n3815 ), .S(st_cfctl) );
    snl_nand14x0 \CODEIF/CNT/U195  ( .ZN(\CODEIF/pgfpoe_in ), .A(
        \CODEIF/CNT/n3793 ), .B(\CODEIF/CNT/n3791 ), .C(\CODEIF/CNT/n3794 ), 
        .D(\CODEIF/CNT/n3795 ) );
    snl_nand03x0 \CODEIF/CNT/U212  ( .ZN(\CODEIF/CNT/n3768 ), .A(
        \CODEIF/CNT/n3809 ), .B(\CODEIF/CNT/n3821 ), .C(\CODEIF/CNT/cst[2] )
         );
    snl_aoi112x0 \CODEIF/CNT/U235  ( .ZN(\CODEIF/CNT/n3792 ), .A(
        \CODEIF/CNT/n3835 ), .B(\CODEIF/CNT/n3797 ), .C(\CODEIF/wprotect0 ), 
        .D(\CODEIF/CNT/n3793 ) );
    snl_aoi012x1 \CODEIF/CNT/U240  ( .ZN(\CODEIF/CNT/n3784 ), .A(
        \CODEIF/CNT/n3827 ), .B(\CODEIF/CNT/n3767 ), .C(\CODEIF/wprotect1 ) );
    snl_invx05 \CODEIF/CNT/U267  ( .ZN(\CODEIF/CNT/n3834 ), .A(
        \CODEIF/CNT/n3825 ) );
    snl_nor02x1 \CODEIF/CNT/U209  ( .ZN(\CODEIF/CNT/n3819 ), .A(
        \CODEIF/CNT/n3801 ), .B(\CODEIF/CNT/cst[3] ) );
    snl_oai122x0 \CODEIF/CNT/U194  ( .ZN(\CODEIF/pgfpce_in ), .A(
        \CODEIF/CNT/n3789 ), .B(\CODEIF/CNT/n3790 ), .C(\CODEIF/CNT/cst[3] ), 
        .D(\CODEIF/CNT/n3791 ), .E(\CODEIF/CNT/n3792 ) );
    snl_ao013x1 \CODEIF/CNT/U200  ( .Z(\CODEIF/CNT/n3806 ), .A(
        \CODEIF/CNT/n3810 ), .B(\CODEIF/CNT/n3809 ), .C(\CODEIF/CNT/n3811 ), 
        .D(\CODEIF/CNT/cst[4] ) );
    snl_ao1b1b3x0 \CODEIF/CNT/U227  ( .Z(\CODEIF/CNT/n3779 ), .A(
        \CODEIF/CNT/n3829 ), .B(\CODEIF/CNT/cst[0] ), .C(\CODEIF/CNT/n3822 ), 
        .D(\CODEIF/CNT/n3830 ), .E(\CODEIF/CNT/n3773 ) );
    snl_invx05 \CODEIF/CNT/U249  ( .ZN(\CODEIF/CNT/n3833 ), .A(
        \CODEIF/CNT/n3826 ) );
    snl_nor03x0 \CODEIF/CNT/U252  ( .ZN(\CODEIF/CNT/n3816 ), .A(
        \CODEIF/CNT/n3821 ), .B(\CODEIF/CNT/n3822 ), .C(\CODEIF/CNT/n3823 ) );
    snl_invx05 \CODEIF/CNT/U275  ( .ZN(\CODEIF/CNT/n3839 ), .A(
        \CODEIF/CNT/n3841 ) );
    snl_ffqrnx1 \CODEIF/CNT/cst_reg[1]  ( .Q(\CODEIF/CNT/cst[1] ), .D(
        \CODEIF/CNT/nst[1] ), .RN(\CODEIF/n3862 ), .CP(SCLK) );
    snl_aoi012x1 \CODEIF/CNT/U201  ( .ZN(\CODEIF/CNT/n3796 ), .A(
        \CODEIF/CNT/n3812 ), .B(\CODEIF/CNT/cst[4] ), .C(\CODEIF/CNT/n3813 )
         );
    snl_invx05 \CODEIF/CNT/U208  ( .ZN(\CODEIF/CNT/n3805 ), .A(
        \CODEIF/CNT/cst[3] ) );
    snl_invx05 \CODEIF/CNT/U213  ( .ZN(\CODEIF/CNT/n3818 ), .A(
        \CODEIF/CNT/cst[4] ) );
    snl_aoi0b12x0 \CODEIF/CNT/U234  ( .ZN(\CODEIF/CNT/n3795 ), .A(
        \CODEIF/CNT/cst[3] ), .B(\CODEIF/CNT/n3797 ), .C(\CODEIF/CNT/n3801 )
         );
    snl_aoi1b12x0 \CODEIF/CNT/U241  ( .ZN(\CODEIF/CNT/n3785 ), .A(cf_wait), 
        .B(\CODEIF/CNT/n3837 ), .C(\CODEIF/CNT/n3781 ), .D(\CODEIF/CNT/n3773 )
         );
    snl_invx05 \CODEIF/CNT/U266  ( .ZN(\CODEIF/CNT/n3838 ), .A(
        \CODEIF/CNT/n3798 ) );
    snl_oai023x0 \CODEIF/CNT/U226  ( .ZN(\CODEIF/CNT/n3773 ), .A(
        \CODEIF/CNT/n3828 ), .B(\CODEIF/CNT/n3821 ), .C(\CODEIF/CNT/n3823 ), 
        .D(\CODEIF/CNT/n3790 ), .E(\CODEIF/CNT/n3799 ) );
    snl_invx05 \CODEIF/CNT/U248  ( .ZN(\CODEIF/CNT/n3803 ), .A(
        \CODEIF/CNT/n3768 ) );
    snl_invx05 \CODEIF/CNT/U253  ( .ZN(\CODEIF/CNT/n3786 ), .A(
        \CODEIF/CNT/n3816 ) );
    snl_nand03x0 \CODEIF/CNT/U274  ( .ZN(\CODEIF/CNT/n3841 ), .A(
        \CODEIF/CNT/n3826 ), .B(\CODEIF/CNT/n3776 ), .C(\CODEIF/CNT/n3777 ) );
    snl_nand02x1 \CODEIF/CNT/U188  ( .ZN(\CODEIF/fddacnt_in ), .A(
        \CODEIF/CNT/n3767 ), .B(\CODEIF/CNT/n3768 ) );
    snl_and02x1 \CODEIF/CNT/U206  ( .Z(\CODEIF/CNT/n3817 ), .A(
        \CODEIF/CNT/n3810 ), .B(\CODEIF/CNT/n3818 ) );
    snl_nor02x1 \CODEIF/CNT/U254  ( .ZN(\CODEIF/CNT/n3807 ), .A(
        \CODEIF/CNT/n3797 ), .B(\CODEIF/CNT/n3814 ) );
    snl_invx05 \CODEIF/CNT/U273  ( .ZN(\CODEIF/CNT/n3837 ), .A(
        \CODEIF/CNT/n3840 ) );
    snl_invx05 \CODEIF/CNT/U268  ( .ZN(\CODEIF/CNT/n3835 ), .A(
        \CODEIF/CNT/n3814 ) );
    snl_nand02x1 \CODEIF/CNT/U214  ( .ZN(\CODEIF/CNT/n3822 ), .A(
        \CODEIF/CNT/cst[4] ), .B(\CODEIF/CNT/n3805 ) );
    snl_nand03x0 \CODEIF/CNT/U221  ( .ZN(\CODEIF/CNT/n3826 ), .A(
        \CODEIF/CNT/n3817 ), .B(\CODEIF/CNT/n3805 ), .C(\CODEIF/CNT/cst[0] )
         );
    snl_aoi012x1 \CODEIF/CNT/U233  ( .ZN(\CODEIF/CNT/n3800 ), .A(
        \CODEIF/CNT/n3833 ), .B(\CODEIF/CNT/n3834 ), .C(\CODEIF/CNT/n3770 ) );
    snl_nand04x0 \CODEIF/CNT/U193  ( .ZN(\CODEIF/CNT/nst[4] ), .A(
        \CODEIF/CNT/n3786 ), .B(\CODEIF/CNT/n3777 ), .C(\CODEIF/CNT/n3787 ), 
        .D(\CODEIF/CNT/n3788 ) );
    snl_nor02x1 \CODEIF/CNT/U246  ( .ZN(\CODEIF/CNT/n3769 ), .A(
        \CODEIF/CNT/n3797 ), .B(\CODEIF/CNT/n3794 ) );
    snl_invx05 \CODEIF/CNT/U261  ( .ZN(\CODEIF/CNT/n3791 ), .A(
        \CODEIF/CNT/n3824 ) );
    snl_aoi123x0 \CODEIF/CNT/U228  ( .ZN(\CODEIF/CNT/n3781 ), .A(
        \CODEIF/CNT/n3827 ), .B(\CODEIF/CNT/n3809 ), .C(\CODEIF/CNT/n3767 ), 
        .D(\CODEIF/CNT/cst[3] ), .E(\CODEIF/CNT/n3824 ), .F(\CODEIF/CNT/n3769 
        ) );
    snl_ao222x1 \REGF/pbmemout1/U8  ( .Z(\pk_adb_h[9] ), .A(\REGF/RO_EACC[9] ), 
        .B(eaccbsel), .C(\REGF/RO_SRDA[9] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[9] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U13  ( .Z(\pk_adb_h[4] ), .A(\REGF/RO_EACC[4] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[4] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[4] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U14  ( .Z(\pk_adb_h[3] ), .A(\REGF/RO_EACC[3] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[3] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[3] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U21  ( .Z(\pk_adb_h[26] ), .A(
        \REGF/RO_EACC[26] ), .B(eaccbsel), .C(\REGF/RO_SRDA[26] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[26] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U54  ( .ZN(\pk_ada_h[10] ), .A(
        \REGF/pbmemout1/n5699 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5700 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U73  ( .ZN(\pk_ada_h[29] ), .A(
        \REGF/pbmemout1/n5737 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5738 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U113  ( .Z(\pk_pdo_h[5] ), .A(
        \REGF/pbmemout1/n5765 ), .B(\REGF/pbmemout1/n5766 ), .C(
        \REGF/pbmemout1/n5767 ), .D(\REGF/pbmemout1/n5768 ) );
    snl_nand04x0 \REGF/pbmemout1/U223  ( .ZN(\REGF/pbmemout1/n5782 ), .A(
        \REGF/pbmemout1/n5888 ), .B(\REGF/pbmemout1/n5887 ), .C(
        \REGF/pbmemout1/n5886 ), .D(\REGF/pbmemout1/n5885 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U432  ( .ZN(\REGF/pbmemout1/n6056 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[28] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[28] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[28] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U840  ( .ZN(\REGF/pbmemout1/n6382 ), .A(
        \REGF/RO_PCON[0] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[0] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[0] ), .F(\pk_rread_h[54] ), .G(
        \pk_stat_h[0] ), .H(\pk_rread_h[55] ) );
    snl_or04x1 \REGF/pbmemout1/U134  ( .Z(\pk_pdo_h[26] ), .A(
        \REGF/pbmemout1/n5849 ), .B(\REGF/pbmemout1/n5850 ), .C(
        \REGF/pbmemout1/n5851 ), .D(\REGF/pbmemout1/n5852 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U692  ( .ZN(\REGF/pbmemout1/n6264 ), .A(
        \pk_s0ba_h[16] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[16] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[16] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[16] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U702  ( .ZN(\REGF/pbmemout1/n6272 ), .A(
        \pk_spr_h[16] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[16] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[16] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[16] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U725  ( .ZN(\REGF/pbmemout1/n6290 ), .A(
        \pk_saseo_h[1] ), .B(\pk_rread_h[4] ), .C(pk_pcser_h), .D(
        \pk_rread_h[5] ), .E(\pk_saco_lh[14] ), .F(\pk_rread_h[6] ), .G(
        \pk_idcz_h[14] ), .H(\pk_rread_h[7] ) );
    snl_oai022x1 \REGF/pbmemout1/U96  ( .ZN(\REGF/pbmemout1/O_LDO[20] ), .A(
        \REGF/pbmemout1/n5719 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5720 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U198  ( .ZN(\REGF/pbmemout1/n5702 ), .A(
        \REGF/RO_EACC[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U204  ( .ZN(\REGF/pbmemout1/n5873 ), .A(
        \pk_rread_h[0] ), .B(1'b0), .C(\pk_rread_h[1] ), .D(1'b0), .E(
        \pk_rread_h[2] ), .F(1'b0), .G(\pk_rread_h[3] ), .H(1'b0) );
    snl_aoi2222x0 \REGF/pbmemout1/U394  ( .ZN(\REGF/pbmemout1/n6025 ), .A(
        \pk_s89l_h[2] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[2] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[2] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[2] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U415  ( .ZN(\REGF/pbmemout1/n6042 ), .A(
        \pk_s01l_h[29] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[29] ), .F(\pk_rread_h[38] ), .G(1'b0), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U585  ( .ZN(\REGF/pbmemout1/n6178 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[20] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[20] ), .H(
        \pk_rread_h[7] ) );
    snl_nand04x0 \REGF/pbmemout1/U338  ( .ZN(\REGF/pbmemout1/n5757 ), .A(
        \REGF/pbmemout1/n5980 ), .B(\REGF/pbmemout1/n5979 ), .C(
        \REGF/pbmemout1/n5978 ), .D(\REGF/pbmemout1/n5977 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U529  ( .ZN(\REGF/pbmemout1/n6133 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U356  ( .ZN(\REGF/pbmemout1/n5995 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[31] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[31] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U371  ( .ZN(\REGF/pbmemout1/n6007 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U560  ( .ZN(\REGF/pbmemout1/n6158 ), .A(
        \REGF/RO_PCON[22] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U619  ( .ZN(\REGF/pbmemout1/n6205 ), .A(
        \REGF/RO_EST2[1] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[1] ), .D(
        \pk_rread_h[49] ), .E(1'b0), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U650  ( .ZN(\REGF/pbmemout1/n6230 ), .A(
        \REGF/pk_s8ba_h[18] ), .B(\pk_rread_h[20] ), .C(\REGF/pk_s7ba_h[18] ), 
        .D(\pk_rread_h[21] ), .E(\REGF/pk_s6ba_h[18] ), .F(\pk_rread_h[22] ), 
        .G(\REGF/pk_s5ba_h[18] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U789  ( .ZN(\REGF/pbmemout1/n6341 ), .A(
        \pk_scba_h[11] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[11] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[11] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[11] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U547  ( .ZN(\REGF/pbmemout1/n6148 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_invx05 \REGF/pbmemout1/U166  ( .ZN(\REGF/pbmemout1/n5732 ), .A(
        \REGF/RO_EACC[26] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U677  ( .ZN(\REGF/pbmemout1/n6252 ), .A(
        \pk_sra1_h[17] ), .B(\pk_rread_h[44] ), .C(CDOUT[17]), .D(
        \pk_rread_h[45] ), .E(CDOUT[49]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[17] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U777  ( .ZN(\REGF/pbmemout1/n6332 ), .A(
        \pk_sra1_h[12] ), .B(\pk_rread_h[44] ), .C(CDOUT[12]), .D(
        \pk_rread_h[45] ), .E(CDOUT[44]), .F(\pk_rread_h[46] ), .G(CDOUT[42]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U809  ( .ZN(\REGF/pbmemout1/n6357 ), .A(
        \pk_scba_h[10] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[10] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[10] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[10] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U256  ( .ZN(\REGF/pbmemout1/n5915 ), .A(
        \REGF/RO_LLPSAS[7] ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[7] ), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[7] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[7] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U447  ( .ZN(\REGF/pbmemout1/n6068 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U271  ( .ZN(\REGF/pbmemout1/n5927 ), .A(
        \pk_s4ba_h[6] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[6] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[6] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[6] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U835  ( .ZN(\REGF/pbmemout1/n6378 ), .A(
        \pk_s01l_h[0] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[0] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[0] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U460  ( .ZN(\REGF/pbmemout1/n6078 ), .A(
        \REGF/RO_PCON[27] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U812  ( .ZN(\REGF/pbmemout1/n6360 ), .A(
        \pk_s0ba_h[10] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[10] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[10] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[10] ), .H(\pk_rread_h[31] ) );
    snl_oai022x1 \REGF/pbmemout1/U68  ( .ZN(\pk_ada_h[24] ), .A(
        \REGF/pbmemout1/n5727 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5728 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U108  ( .Z(\pk_pdo_h[0] ), .A(
        \REGF/pbmemout1/n5745 ), .B(\REGF/pbmemout1/n5746 ), .C(
        \REGF/pbmemout1/n5747 ), .D(\REGF/pbmemout1/n5748 ) );
    snl_invx05 \REGF/pbmemout1/U141  ( .ZN(\REGF/pbmemout1/n5697 ), .A(
        \REGF/RO_ACC[9] ) );
    snl_invx05 \REGF/pbmemout1/U183  ( .ZN(\REGF/pbmemout1/n5717 ), .A(
        \REGF/RO_ACC[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U294  ( .ZN(\REGF/pbmemout1/n5945 ), .A(
        \pk_s89l_h[5] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[5] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[5] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[5] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U304  ( .ZN(\REGF/pbmemout1/n5953 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(
        \REGF/pk_scti_h[4] ), .F(\pk_rread_h[2] ), .G(1'b0), .H(
        \pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U485  ( .ZN(\REGF/pbmemout1/n6098 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(1'b0), .F(
        \pk_rread_h[6] ), .G(\REGF/pk_idcz_h[25] ), .H(\pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U750  ( .ZN(\REGF/pbmemout1/n6310 ), .A(
        \pk_s8ba_h[13] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[13] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[13] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[13] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U515  ( .ZN(\REGF/pbmemout1/n6122 ), .A(
        \pk_s01l_h[24] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[20] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[24] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U625  ( .ZN(\REGF/pbmemout1/n6210 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[19] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[19] ), .H(
        \pk_rread_h[7] ) );
    snl_nand04x0 \REGF/pbmemout1/U323  ( .ZN(\REGF/pbmemout1/n5762 ), .A(
        \REGF/pbmemout1/n5968 ), .B(\REGF/pbmemout1/n5967 ), .C(
        \REGF/pbmemout1/n5966 ), .D(\REGF/pbmemout1/n5965 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U532  ( .ZN(\REGF/pbmemout1/n6136 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[23] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[23] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[23] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U602  ( .ZN(\REGF/pbmemout1/n6192 ), .A(
        \pk_spr_h[20] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[20] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[20] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[20] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U792  ( .ZN(\REGF/pbmemout1/n6344 ), .A(
        \pk_s0ba_h[11] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[11] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[11] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[11] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U238  ( .ZN(\REGF/pbmemout1/n5777 ), .A(
        \REGF/pbmemout1/n5900 ), .B(\REGF/pbmemout1/n5899 ), .C(
        \REGF/pbmemout1/n5898 ), .D(\REGF/pbmemout1/n5897 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U689  ( .ZN(\REGF/pbmemout1/n6261 ), .A(
        \pk_scba_h[16] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[16] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[16] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[16] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U719  ( .ZN(\REGF/pbmemout1/n6285 ), .A(
        \REGF/RO_EST2[15] ), .B(\pk_rread_h[48] ), .C(ph_tirtendh), .D(
        \pk_rread_h[49] ), .E(1'b0), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U429  ( .ZN(\REGF/pbmemout1/n6053 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_invx05 \REGF/pbmemout1/U174  ( .ZN(\REGF/pbmemout1/n5724 ), .A(
        \REGF/RO_EACC[22] ) );
    snl_invx05 \REGF/pbmemout1/U191  ( .ZN(\REGF/pbmemout1/n5709 ), .A(
        \REGF/RO_ACC[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U286  ( .ZN(\REGF/pbmemout1/n5939 ), .A(
        \pk_idcy_h[5] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[5] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[5] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[5] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U507  ( .ZN(\REGF/pbmemout1/n6116 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U316  ( .ZN(\REGF/pbmemout1/n5963 ), .A(
        \REGF/RO_LLPSAS[4] ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[4] ), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[4] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[4] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U497  ( .ZN(\REGF/pbmemout1/n6108 ), .A(1'b0
        ), .B(\pk_rread_h[44] ), .C(CDOUT[25]), .D(\pk_rread_h[45] ), .E(CDOUT
        [57]), .F(\pk_rread_h[46] ), .G(\REGF/RO_DDCS[25] ), .H(
        \pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U637  ( .ZN(\REGF/pbmemout1/n6220 ), .A(
        \pk_sra1_h[19] ), .B(\pk_rread_h[44] ), .C(CDOUT[19]), .D(
        \pk_rread_h[45] ), .E(CDOUT[51]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[19] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U780  ( .ZN(\REGF/pbmemout1/n6334 ), .A(
        \REGF/RO_PCON[12] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[12] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[12] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U331  ( .ZN(\REGF/pbmemout1/n5975 ), .A(
        \pk_s4ba_h[3] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[3] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[3] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[3] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U610  ( .ZN(\REGF/pbmemout1/n6198 ), .A(
        \pk_s8ba_h[1] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[1] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[1] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[1] ), .H(\pk_rread_h[23] ) );
    snl_nand04x0 \REGF/pbmemout1/U378  ( .ZN(\REGF/pbmemout1/n5865 ), .A(
        \REGF/pbmemout1/n6012 ), .B(\REGF/pbmemout1/n6011 ), .C(
        \REGF/pbmemout1/n6010 ), .D(\REGF/pbmemout1/n6009 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U520  ( .ZN(\REGF/pbmemout1/n6126 ), .A(
        \REGF/RO_PCON[24] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U569  ( .ZN(\REGF/pbmemout1/n6165 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U659  ( .ZN(\REGF/pbmemout1/n6237 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[18] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U244  ( .ZN(\REGF/pbmemout1/n5905 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(
        \REGF/pk_scti_h[7] ), .F(\pk_rread_h[2] ), .G(1'b0), .H(
        \pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U765  ( .ZN(\REGF/pbmemout1/n6322 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[12] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[12] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U827  ( .ZN(\REGF/pbmemout1/n6372 ), .A(
        \pk_pcs1_h[0] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[0] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[0] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[0] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U455  ( .ZN(\REGF/pbmemout1/n6074 ), .A(
        \pk_s01l_h[27] ), .B(\pk_rread_h[36] ), .C(\REGF/RO_TRCO[27] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[27] ), .H(\pk_rread_h[39] ) );
    snl_ao222x1 \REGF/pbmemout1/U28  ( .Z(\pk_adb_h[1] ), .A(\REGF/RO_EACC[1] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[1] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[1] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U33  ( .Z(\pk_adb_h[15] ), .A(
        \REGF/RO_EACC[15] ), .B(eaccbsel), .C(\REGF/RO_SRDA[15] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[15] ), .F(accbsel) );
    snl_nand04x0 \REGF/pbmemout1/U263  ( .ZN(\REGF/pbmemout1/n5774 ), .A(
        \REGF/pbmemout1/n5920 ), .B(\REGF/pbmemout1/n5919 ), .C(
        \REGF/pbmemout1/n5918 ), .D(\REGF/pbmemout1/n5917 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U472  ( .ZN(\REGF/pbmemout1/n6088 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[26] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[26] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[26] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U800  ( .ZN(\REGF/pbmemout1/n6350 ), .A(
        \REGF/RO_PCON[11] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[11] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[11] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_invx05 \REGF/pbmemout1/U148  ( .ZN(\REGF/pbmemout1/n5690 ), .A(
        \REGF/RO_EACC[5] ) );
    snl_invx05 \REGF/pbmemout1/U153  ( .ZN(\REGF/pbmemout1/n5685 ), .A(
        \REGF/RO_ACC[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U742  ( .ZN(\REGF/pbmemout1/n6304 ), .A(
        \pk_spr_h[14] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[14] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[14] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[14] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U759  ( .ZN(\REGF/pbmemout1/n6317 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[43]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_ao222x1 \REGF/pbmemout1/U34  ( .Z(\pk_adb_h[14] ), .A(
        \REGF/RO_EACC[14] ), .B(eaccbsel), .C(\REGF/RO_SRDA[14] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[14] ), .F(accbsel) );
    snl_invx1 \REGF/pbmemout1/U41  ( .ZN(\REGF/pbmemout1/n5680 ), .A(eaccasel)
         );
    snl_oai022x1 \REGF/pbmemout1/U46  ( .ZN(\pk_ada_h[2] ), .A(
        \REGF/pbmemout1/n5683 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5684 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U61  ( .ZN(\pk_ada_h[17] ), .A(
        \REGF/pbmemout1/n5713 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5714 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U84  ( .ZN(\REGF/pbmemout1/O_LDO[8] ), .A(
        \REGF/pbmemout1/n5695 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5696 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_nand04x0 \REGF/pbmemout1/U278  ( .ZN(\REGF/pbmemout1/n5769 ), .A(
        \REGF/pbmemout1/n5932 ), .B(\REGF/pbmemout1/n5931 ), .C(
        \REGF/pbmemout1/n5930 ), .D(\REGF/pbmemout1/n5929 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U469  ( .ZN(\REGF/pbmemout1/n6085 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U344  ( .ZN(\REGF/pbmemout1/n5985 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U363  ( .ZN(\REGF/pbmemout1/n5870 ), .A(
        \REGF/pbmemout1/n6000 ), .B(\REGF/pbmemout1/n5999 ), .C(
        \REGF/pbmemout1/n5998 ), .D(\REGF/pbmemout1/n5997 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U642  ( .ZN(\REGF/pbmemout1/n6224 ), .A(
        \pk_spr_h[19] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[19] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[19] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[19] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U555  ( .ZN(\REGF/pbmemout1/n6154 ), .A(
        \pk_s01l_h[22] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[18] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[22] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[22] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U572  ( .ZN(\REGF/pbmemout1/n6168 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[21] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[21] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[21] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U665  ( .ZN(\REGF/pbmemout1/n6242 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[17] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[17] ), .H(
        \pk_rread_h[7] ) );
    snl_oai022x1 \REGF/pbmemout1/U101  ( .ZN(\REGF/pbmemout1/O_LDO[25] ), .A(
        \REGF/pbmemout1/n5729 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5730 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U231  ( .ZN(\REGF/pbmemout1/n5895 ), .A(
        \pk_s4ba_h[8] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[8] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[8] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[8] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U420  ( .ZN(\REGF/pbmemout1/n6046 ), .A(
        \REGF/RO_PCON[29] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U710  ( .ZN(\REGF/pbmemout1/n6278 ), .A(
        \pk_s8ba_h[15] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[15] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[15] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[15] ), .H(\pk_rread_h[23] ) );
    snl_or04x1 \REGF/pbmemout1/U126  ( .Z(\pk_pdo_h[18] ), .A(
        \REGF/pbmemout1/n5817 ), .B(\REGF/pbmemout1/n5818 ), .C(
        \REGF/pbmemout1/n5819 ), .D(\REGF/pbmemout1/n5820 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U680  ( .ZN(\REGF/pbmemout1/n6254 ), .A(
        \REGF/RO_PCON[17] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[17] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[17] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U737  ( .ZN(\REGF/pbmemout1/n6300 ), .A(
        \pk_sra1_h[14] ), .B(\pk_rread_h[44] ), .C(CDOUT[14]), .D(
        \pk_rread_h[45] ), .E(CDOUT[46]), .F(\pk_rread_h[46] ), .G(CDOUT[44]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U211  ( .ZN(\REGF/pbmemout1/n5879 ), .A(
        \pk_rread_h[24] ), .B(\pk_s4ba_h[9] ), .C(\pk_rread_h[25] ), .D(
        \pk_s3ba_h[9] ), .E(\pk_rread_h[26] ), .F(\pk_s2ba_h[9] ), .G(
        \pk_rread_h[27] ), .H(\pk_s1ba_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U216  ( .ZN(\REGF/pbmemout1/n5883 ), .A(
        \pk_rread_h[40] ), .B(\REGF/RO_LLPSAS[9] ), .C(\pk_rread_h[41] ), .D(
        1'b0), .E(\pk_rread_h[42] ), .F(\REGF/RO_SRDA[9] ), .G(
        \pk_rread_h[43] ), .H(\pk_sra2_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U597  ( .ZN(\REGF/pbmemout1/n6188 ), .A(
        \pk_sra1_h[20] ), .B(\pk_rread_h[44] ), .C(CDOUT[20]), .D(
        \pk_rread_h[45] ), .E(CDOUT[52]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[20] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U381  ( .ZN(\REGF/pbmemout1/n6015 ), .A(
        \REGF/pk_indz_h[30] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[30] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[30] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[30] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U386  ( .ZN(\REGF/pbmemout1/n6019 ), .A(
        \pk_idcy_h[2] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[2] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[2] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[2] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U407  ( .ZN(\REGF/pbmemout1/n6036 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U400  ( .ZN(\REGF/pbmemout1/n6030 ), .A(
        \REGF/RO_PCON[2] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[2] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[2] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U590  ( .ZN(\REGF/pbmemout1/n6182 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_oai022x1 \REGF/pbmemout1/U66  ( .ZN(\pk_ada_h[22] ), .A(
        \REGF/pbmemout1/n5723 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5724 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U106  ( .ZN(\REGF/pbmemout1/O_LDO[30] ), .A(
        \REGF/pbmemout1/n5739 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5740 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U121  ( .Z(\pk_pdo_h[13] ), .A(
        \REGF/pbmemout1/n5797 ), .B(\REGF/pbmemout1/n5798 ), .C(
        \REGF/pbmemout1/n5799 ), .D(\REGF/pbmemout1/n5800 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U730  ( .ZN(\REGF/pbmemout1/n6294 ), .A(
        \pk_s8ba_h[14] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[14] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[14] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[14] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U687  ( .ZN(\REGF/pbmemout1/n6260 ), .A(
        \pk_pcs1_h[16] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[16] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[16] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[16] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U236  ( .ZN(\REGF/pbmemout1/n5899 ), .A(
        \REGF/RO_LLPSAS[8] ), .B(\pk_rread_h[40] ), .C(1'b0), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[8] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[8] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U717  ( .ZN(\REGF/pbmemout1/n6284 ), .A(
        \pk_sra1_h[15] ), .B(\pk_rread_h[44] ), .C(CDOUT[15]), .D(
        \pk_rread_h[45] ), .E(CDOUT[47]), .F(\pk_rread_h[46] ), .G(1'b0), .H(
        \pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U427  ( .ZN(\REGF/pbmemout1/n6052 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_oai022x1 \REGF/pbmemout1/U83  ( .ZN(\REGF/pbmemout1/O_LDO[7] ), .A(
        \REGF/pbmemout1/n5693 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5694 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U168  ( .ZN(\REGF/pbmemout1/n5730 ), .A(
        \REGF/RO_EACC[25] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U779  ( .ZN(\REGF/pbmemout1/n6333 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[42]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U258  ( .ZN(\REGF/pbmemout1/n5773 ), .A(
        \REGF/pbmemout1/n5916 ), .B(\REGF/pbmemout1/n5915 ), .C(
        \REGF/pbmemout1/n5914 ), .D(\REGF/pbmemout1/n5913 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U449  ( .ZN(\REGF/pbmemout1/n6069 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U662  ( .ZN(\REGF/pbmemout1/n6240 ), .A(
        \pk_spr_h[18] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[18] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[18] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[18] ), .H(\pk_rread_h[63] ) );
    snl_oai022x1 \REGF/pbmemout1/U98  ( .ZN(\REGF/pbmemout1/O_LDO[22] ), .A(
        \REGF/pbmemout1/n5723 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5724 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_nand04x0 \REGF/pbmemout1/U343  ( .ZN(\REGF/pbmemout1/n5758 ), .A(
        \REGF/pbmemout1/n5984 ), .B(\REGF/pbmemout1/n5983 ), .C(
        \REGF/pbmemout1/n5982 ), .D(\REGF/pbmemout1/n5981 ) );
    snl_nand04x0 \REGF/pbmemout1/U358  ( .ZN(\REGF/pbmemout1/n5869 ), .A(
        \REGF/pbmemout1/n5996 ), .B(\REGF/pbmemout1/n5995 ), .C(
        \REGF/pbmemout1/n5994 ), .D(\REGF/pbmemout1/n5993 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U364  ( .ZN(\REGF/pbmemout1/n6001 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U552  ( .ZN(\REGF/pbmemout1/n6152 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[22] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[22] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[22] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U575  ( .ZN(\REGF/pbmemout1/n6170 ), .A(
        \pk_s01l_h[21] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[17] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[21] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[21] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U645  ( .ZN(\REGF/pbmemout1/n6226 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[18] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[18] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U549  ( .ZN(\REGF/pbmemout1/n6149 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_invx05 \REGF/pbmemout1/U154  ( .ZN(\REGF/pbmemout1/n5742 ), .A(
        \REGF/RO_EACC[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U679  ( .ZN(\REGF/pbmemout1/n6253 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[17] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U745  ( .ZN(\REGF/pbmemout1/n6306 ), .A(
        \pk_saseo_h[0] ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), 
        .E(\pk_saco_lh[13] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[13] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U264  ( .ZN(\REGF/pbmemout1/n5921 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(
        \REGF/pk_scti_h[6] ), .F(\pk_rread_h[2] ), .G(1'b0), .H(
        \pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U475  ( .ZN(\REGF/pbmemout1/n6090 ), .A(
        \pk_s01l_h[26] ), .B(\pk_rread_h[36] ), .C(\REGF/RO_TRCO[26] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[26] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U807  ( .ZN(\REGF/pbmemout1/n6356 ), .A(
        \pk_pcs1_h[10] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[10] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[10] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[10] ), .H(\pk_rread_h[15] ) );
    snl_ao222x1 \REGF/pbmemout1/U26  ( .Z(\pk_adb_h[21] ), .A(
        \REGF/RO_EACC[21] ), .B(eaccbsel), .C(\REGF/RO_SRDA[21] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[21] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U48  ( .ZN(\pk_ada_h[4] ), .A(
        \REGF/pbmemout1/n5687 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5688 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U128  ( .Z(\pk_pdo_h[20] ), .A(
        \REGF/pbmemout1/n5825 ), .B(\REGF/pbmemout1/n5826 ), .C(
        \REGF/pbmemout1/n5827 ), .D(\REGF/pbmemout1/n5828 ) );
    snl_invx05 \REGF/pbmemout1/U173  ( .ZN(\REGF/pbmemout1/n5725 ), .A(
        \REGF/RO_ACC[23] ) );
    snl_nand04x0 \REGF/pbmemout1/U243  ( .ZN(\REGF/pbmemout1/n5778 ), .A(
        \REGF/pbmemout1/n5904 ), .B(\REGF/pbmemout1/n5903 ), .C(
        \REGF/pbmemout1/n5902 ), .D(\REGF/pbmemout1/n5901 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U452  ( .ZN(\REGF/pbmemout1/n6072 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[27] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[27] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[27] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U762  ( .ZN(\REGF/pbmemout1/n6320 ), .A(
        \pk_spr_h[13] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[13] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[13] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[13] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U820  ( .ZN(\REGF/pbmemout1/n6366 ), .A(
        \REGF/RO_PCON[10] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[10] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[10] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_invx05 \REGF/pbmemout1/U184  ( .ZN(\REGF/pbmemout1/n5716 ), .A(
        \REGF/RO_EACC[18] ) );
    snl_invx05 \REGF/pbmemout1/U196  ( .ZN(\REGF/pbmemout1/n5704 ), .A(
        \REGF/RO_EACC[12] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U336  ( .ZN(\REGF/pbmemout1/n5979 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[3] ), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[3] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[3] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U527  ( .ZN(\REGF/pbmemout1/n6132 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U617  ( .ZN(\REGF/pbmemout1/n6204 ), .A(
        \pk_sra1_h[1] ), .B(\pk_rread_h[44] ), .C(CDOUT[1]), .D(
        \pk_rread_h[45] ), .E(CDOUT[33]), .F(\pk_rread_h[46] ), .G(1'b0), .H(
        \pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U281  ( .ZN(\REGF/pbmemout1/n5935 ), .A(
        \pk_indz_h[6] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[6] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[6] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[6] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U311  ( .ZN(\REGF/pbmemout1/n5959 ), .A(
        \pk_s4ba_h[4] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[4] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[4] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[4] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U630  ( .ZN(\REGF/pbmemout1/n6214 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U787  ( .ZN(\REGF/pbmemout1/n6340 ), .A(
        \pk_pcs1_h[11] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[11] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[11] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[11] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U490  ( .ZN(\REGF/pbmemout1/n6102 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U324  ( .ZN(\REGF/pbmemout1/n5969 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(\REGF/pk_exco_h[3] ), .D(\pk_rread_h[1] ), 
        .E(\REGF/pk_scti_h[3] ), .F(\pk_rread_h[2] ), .G(1'b0), .H(
        \pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U500  ( .ZN(\REGF/pbmemout1/n6110 ), .A(
        \REGF/RO_PCON[25] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U535  ( .ZN(\REGF/pbmemout1/n6138 ), .A(
        \pk_s01l_h[23] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[19] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[23] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[23] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U605  ( .ZN(\REGF/pbmemout1/n6194 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[1] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[1] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U795  ( .ZN(\REGF/pbmemout1/n6346 ), .A(
        \pk_s01l_h[11] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[11] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[11] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[11] ), .H(\pk_rread_h[39] ) );
    snl_nand04x0 \REGF/pbmemout1/U293  ( .ZN(\REGF/pbmemout1/n5768 ), .A(
        \REGF/pbmemout1/n5944 ), .B(\REGF/pbmemout1/n5943 ), .C(
        \REGF/pbmemout1/n5942 ), .D(\REGF/pbmemout1/n5941 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U622  ( .ZN(\REGF/pbmemout1/n6208 ), .A(
        \pk_spr_h[1] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[1] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[1] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[1] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U303  ( .ZN(\REGF/pbmemout1/n5766 ), .A(
        \REGF/pbmemout1/n5952 ), .B(\REGF/pbmemout1/n5951 ), .C(
        \REGF/pbmemout1/n5950 ), .D(\REGF/pbmemout1/n5949 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U512  ( .ZN(\REGF/pbmemout1/n6120 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[24] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[24] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[24] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U482  ( .ZN(\REGF/pbmemout1/n6096 ), .A(1'b0
        ), .B(\pk_rread_h[60] ), .C(1'b0), .D(\pk_rread_h[61] ), .E(
        \REGF/RO_EACC[26] ), .F(\pk_rread_h[62] ), .G(\REGF/RO_ACC[26] ), .H(
        \pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U739  ( .ZN(\REGF/pbmemout1/n6301 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(ph_byrtendh), .D(\pk_rread_h[49] ), .E(
        CDOUT[44]), .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_invx05 \REGF/pbmemout1/U146  ( .ZN(\REGF/pbmemout1/n5692 ), .A(
        \REGF/RO_EACC[6] ) );
    snl_nand04x0 \REGF/pbmemout1/U218  ( .ZN(\REGF/pbmemout1/n5781 ), .A(
        \REGF/pbmemout1/n5884 ), .B(\REGF/pbmemout1/n5883 ), .C(
        \REGF/pbmemout1/n5882 ), .D(\REGF/pbmemout1/n5881 ) );
    snl_nand04x0 \REGF/pbmemout1/U388  ( .ZN(\REGF/pbmemout1/n5755 ), .A(
        \REGF/pbmemout1/n6020 ), .B(\REGF/pbmemout1/n6019 ), .C(
        \REGF/pbmemout1/n6018 ), .D(\REGF/pbmemout1/n6017 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U599  ( .ZN(\REGF/pbmemout1/n6189 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[20] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U409  ( .ZN(\REGF/pbmemout1/n6037 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U757  ( .ZN(\REGF/pbmemout1/n6316 ), .A(
        \pk_sra1_h[13] ), .B(\pk_rread_h[44] ), .C(CDOUT[13]), .D(
        \pk_rread_h[45] ), .E(CDOUT[45]), .F(\pk_rread_h[46] ), .G(CDOUT[43]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U251  ( .ZN(\REGF/pbmemout1/n5911 ), .A(
        \pk_s4ba_h[7] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[7] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[7] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[7] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U276  ( .ZN(\REGF/pbmemout1/n5931 ), .A(
        \REGF/RO_LLPSAS[6] ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[6] ), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[6] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[6] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U467  ( .ZN(\REGF/pbmemout1/n6084 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U815  ( .ZN(\REGF/pbmemout1/n6362 ), .A(
        \pk_s01l_h[10] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[10] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[10] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[10] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U832  ( .ZN(\REGF/pbmemout1/n6376 ), .A(
        \pk_s0ba_h[0] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[0] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[0] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[0] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U440  ( .ZN(\REGF/pbmemout1/n6062 ), .A(
        \REGF/RO_PCON[28] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_ao222x1 \REGF/pbmemout1/U9  ( .Z(\pk_adb_h[8] ), .A(\REGF/RO_EACC[8] ), 
        .B(eaccbsel), .C(\REGF/RO_SRDA[8] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[8] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U12  ( .Z(\pk_adb_h[5] ), .A(\REGF/RO_EACC[5] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[5] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[5] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U35  ( .Z(\pk_adb_h[13] ), .A(
        \REGF/RO_EACC[13] ), .B(eaccbsel), .C(\REGF/RO_SRDA[13] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[13] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U53  ( .ZN(\pk_ada_h[9] ), .A(
        \REGF/pbmemout1/n5697 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5698 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U91  ( .ZN(\REGF/pbmemout1/O_LDO[15] ), .A(
        \REGF/pbmemout1/n5709 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5710 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U161  ( .ZN(\REGF/pbmemout1/n5737 ), .A(
        \REGF/RO_ACC[29] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U670  ( .ZN(\REGF/pbmemout1/n6246 ), .A(
        \pk_s8ba_h[17] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[17] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[17] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[17] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U770  ( .ZN(\REGF/pbmemout1/n6326 ), .A(
        \pk_s8ba_h[12] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[12] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[12] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[12] ), .H(\pk_rread_h[23] ) );
    snl_invx05 \REGF/pbmemout1/U203  ( .ZN(\REGF/pbmemout1/n5677 ), .A(
        \REGF/RO_ACC[0] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U351  ( .ZN(\REGF/pbmemout1/n5991 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U540  ( .ZN(\REGF/pbmemout1/n6142 ), .A(
        \REGF/RO_PCON[23] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U376  ( .ZN(\REGF/pbmemout1/n6011 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[30] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[30] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U567  ( .ZN(\REGF/pbmemout1/n6164 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U657  ( .ZN(\REGF/pbmemout1/n6236 ), .A(
        \pk_sra1_h[18] ), .B(\pk_rread_h[44] ), .C(CDOUT[18]), .D(
        \pk_rread_h[45] ), .E(CDOUT[50]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[18] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U829  ( .ZN(\REGF/pbmemout1/n6373 ), .A(
        \pk_scba_h[0] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[0] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[0] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[0] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U393  ( .ZN(\REGF/pbmemout1/n5756 ), .A(
        \REGF/pbmemout1/n6024 ), .B(\REGF/pbmemout1/n6023 ), .C(
        \REGF/pbmemout1/n6022 ), .D(\REGF/pbmemout1/n6021 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U582  ( .ZN(\REGF/pbmemout1/n6176 ), .A(
        \pk_spr_h[21] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[21] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[21] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[21] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U412  ( .ZN(\REGF/pbmemout1/n6040 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[29] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[29] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[29] ), .H(
        \pk_rread_h[31] ) );
    snl_oai022x1 \REGF/pbmemout1/U74  ( .ZN(\pk_ada_h[30] ), .A(
        \REGF/pbmemout1/n5739 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5740 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U114  ( .Z(\pk_pdo_h[6] ), .A(
        \REGF/pbmemout1/n5769 ), .B(\REGF/pbmemout1/n5770 ), .C(
        \REGF/pbmemout1/n5771 ), .D(\REGF/pbmemout1/n5772 ) );
    snl_or04x1 \REGF/pbmemout1/U133  ( .Z(\pk_pdo_h[25] ), .A(
        \REGF/pbmemout1/n5845 ), .B(\REGF/pbmemout1/n5846 ), .C(
        \REGF/pbmemout1/n5847 ), .D(\REGF/pbmemout1/n5848 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U695  ( .ZN(\REGF/pbmemout1/n6266 ), .A(
        \pk_s01l_h[16] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[12] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[16] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[16] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U705  ( .ZN(\REGF/pbmemout1/n6274 ), .A(
        pk_sasea_h), .B(\pk_rread_h[4] ), .C(pk_pcsee_h), .D(\pk_rread_h[5] ), 
        .E(\pk_saco_lh[15] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[15] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U722  ( .ZN(\REGF/pbmemout1/n6288 ), .A(
        \pk_spr_h[15] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[15] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[15] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[15] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U224  ( .ZN(\REGF/pbmemout1/n5889 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U435  ( .ZN(\REGF/pbmemout1/n6058 ), .A(
        \pk_s01l_h[28] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[28] ), .F(\pk_rread_h[38] ), .G(1'b0), .H(
        \pk_rread_h[39] ) );
    snl_oai022x1 \REGF/pbmemout1/U99  ( .ZN(\REGF/pbmemout1/O_LDO[23] ), .A(
        \REGF/pbmemout1/n5725 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5726 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U197  ( .ZN(\REGF/pbmemout1/n5703 ), .A(
        \REGF/RO_ACC[12] ) );
    snl_nand04x0 \REGF/pbmemout1/U288  ( .ZN(\REGF/pbmemout1/n5767 ), .A(
        \REGF/pbmemout1/n5940 ), .B(\REGF/pbmemout1/n5939 ), .C(
        \REGF/pbmemout1/n5938 ), .D(\REGF/pbmemout1/n5937 ) );
    snl_nand04x0 \REGF/pbmemout1/U318  ( .ZN(\REGF/pbmemout1/n5761 ), .A(
        \REGF/pbmemout1/n5964 ), .B(\REGF/pbmemout1/n5963 ), .C(
        \REGF/pbmemout1/n5962 ), .D(\REGF/pbmemout1/n5961 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U509  ( .ZN(\REGF/pbmemout1/n6117 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U337  ( .ZN(\REGF/pbmemout1/n5980 ), .A(
        \pk_sra1_h[3] ), .B(\pk_rread_h[44] ), .C(CDOUT[3]), .D(
        \pk_rread_h[45] ), .E(CDOUT[35]), .F(\pk_rread_h[46] ), .G(CDOUT[33]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U499  ( .ZN(\REGF/pbmemout1/n6109 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_DDCS[25] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U639  ( .ZN(\REGF/pbmemout1/n6221 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[19] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U526  ( .ZN(\REGF/pbmemout1/n6131 ), .A(
        \pk_idcy_h[23] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[23] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[23] ), .F(\pk_rread_h[10] ), .G(1'b0), 
        .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U786  ( .ZN(\REGF/pbmemout1/n6339 ), .A(
        \pk_idcy_h[11] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[11] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[11] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[11] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U280  ( .ZN(\REGF/pbmemout1/n5934 ), .A(
        \REGF/RO_PCON[6] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[6] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[6] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U501  ( .ZN(\REGF/pbmemout1/n6111 ), .A(
        \REGF/pk_indz_h[25] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[25] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[25] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[25] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U616  ( .ZN(\REGF/pbmemout1/n6203 ), .A(
        \REGF/RO_LLPSAS[1] ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[1] ), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[1] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[1] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U631  ( .ZN(\REGF/pbmemout1/n6215 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U310  ( .ZN(\REGF/pbmemout1/n5958 ), .A(
        \pk_s8ba_h[4] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[4] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[4] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[4] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U491  ( .ZN(\REGF/pbmemout1/n6103 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_invx05 \REGF/pbmemout1/U155  ( .ZN(\REGF/pbmemout1/n5741 ), .A(
        pk_sign_h) );
    snl_aoi2222x0 \REGF/pbmemout1/U359  ( .ZN(\REGF/pbmemout1/n5997 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[59]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U548  ( .ZN(\REGF/pbmemout1/n5835 ), .A(
        \REGF/pbmemout1/n6148 ), .B(\REGF/pbmemout1/n6147 ), .C(
        \REGF/pbmemout1/n6146 ), .D(\REGF/pbmemout1/n6145 ) );
    snl_nand04x0 \REGF/pbmemout1/U678  ( .ZN(\REGF/pbmemout1/n5813 ), .A(
        \REGF/pbmemout1/n6252 ), .B(\REGF/pbmemout1/n6251 ), .C(
        \REGF/pbmemout1/n6250 ), .D(\REGF/pbmemout1/n6249 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U744  ( .ZN(\REGF/pbmemout1/n6305 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U265  ( .ZN(\REGF/pbmemout1/n5922 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[6] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[6] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U474  ( .ZN(\REGF/pbmemout1/n6089 ), .A(
        \pk_s89l_h[26] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[26] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[26] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[26] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U806  ( .ZN(\REGF/pbmemout1/n6355 ), .A(
        \pk_idcy_h[10] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[10] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[10] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[10] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U242  ( .ZN(\REGF/pbmemout1/n5904 ), .A(
        \pk_spr_h[8] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[8] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[8] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[8] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U453  ( .ZN(\REGF/pbmemout1/n5856 ), .A(
        \REGF/pbmemout1/n6072 ), .B(\REGF/pbmemout1/n6071 ), .C(
        \REGF/pbmemout1/n6070 ), .D(\REGF/pbmemout1/n6069 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U821  ( .ZN(\REGF/pbmemout1/n6367 ), .A(
        \pk_indz_h[10] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[10] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[10] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[10] ), .H(\pk_rread_h[59] ) );
    snl_ao222x1 \REGF/pbmemout1/U27  ( .Z(\pk_adb_h[20] ), .A(
        \REGF/RO_EACC[20] ), .B(eaccbsel), .C(\REGF/RO_SRDA[20] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[20] ), .F(accbsel) );
    snl_invx1 \REGF/pbmemout1/U40  ( .ZN(\REGF/pbmemout1/n5743 ), .A(
        po_raccl_h) );
    snl_oai022x1 \REGF/pbmemout1/U82  ( .ZN(\REGF/pbmemout1/O_LDO[6] ), .A(
        \REGF/pbmemout1/n5691 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5692 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U169  ( .ZN(\REGF/pbmemout1/n5729 ), .A(
        \REGF/RO_ACC[25] ) );
    snl_invx05 \REGF/pbmemout1/U172  ( .ZN(\REGF/pbmemout1/n5726 ), .A(
        \REGF/RO_EACC[23] ) );
    snl_nand04x0 \REGF/pbmemout1/U763  ( .ZN(\REGF/pbmemout1/n5798 ), .A(
        \REGF/pbmemout1/n6320 ), .B(\REGF/pbmemout1/n6319 ), .C(
        \REGF/pbmemout1/n6318 ), .D(\REGF/pbmemout1/n6317 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U259  ( .ZN(\REGF/pbmemout1/n5917 ), .A(
        \REGF/RO_PSTA[20] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[7] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[37]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U778  ( .ZN(\REGF/pbmemout1/n5793 ), .A(
        \REGF/pbmemout1/n6332 ), .B(\REGF/pbmemout1/n6331 ), .C(
        \REGF/pbmemout1/n6330 ), .D(\REGF/pbmemout1/n6329 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U342  ( .ZN(\REGF/pbmemout1/n5984 ), .A(
        \pk_spr_h[3] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[3] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[3] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[3] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U448  ( .ZN(\REGF/pbmemout1/n5855 ), .A(
        \REGF/pbmemout1/n6068 ), .B(\REGF/pbmemout1/n6067 ), .C(
        \REGF/pbmemout1/n6066 ), .D(\REGF/pbmemout1/n6065 ) );
    snl_nand04x0 \REGF/pbmemout1/U553  ( .ZN(\REGF/pbmemout1/n5836 ), .A(
        \REGF/pbmemout1/n6152 ), .B(\REGF/pbmemout1/n6151 ), .C(
        \REGF/pbmemout1/n6150 ), .D(\REGF/pbmemout1/n6149 ) );
    snl_nand04x0 \REGF/pbmemout1/U663  ( .ZN(\REGF/pbmemout1/n5818 ), .A(
        \REGF/pbmemout1/n6240 ), .B(\REGF/pbmemout1/n6239 ), .C(
        \REGF/pbmemout1/n6238 ), .D(\REGF/pbmemout1/n6237 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U365  ( .ZN(\REGF/pbmemout1/n6002 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_hh[30] ), .F(\pk_rread_h[6] ), .G(\REGF/pk_idcz_h[30] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U574  ( .ZN(\REGF/pbmemout1/n6169 ), .A(
        \pk_s89l_h[21] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[21] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[21] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[21] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U644  ( .ZN(\REGF/pbmemout1/n6225 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_oai022x1 \REGF/pbmemout1/U52  ( .ZN(\pk_ada_h[8] ), .A(
        \REGF/pbmemout1/n5695 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5696 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U67  ( .ZN(\pk_ada_h[23] ), .A(
        \REGF/pbmemout1/n5725 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5726 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U107  ( .ZN(\REGF/pbmemout1/O_LDO[31] ), .A(
        \REGF/pbmemout1/n5741 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5742 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U120  ( .Z(\pk_pdo_h[12] ), .A(
        \REGF/pbmemout1/n5793 ), .B(\REGF/pbmemout1/n5794 ), .C(
        \REGF/pbmemout1/n5795 ), .D(\REGF/pbmemout1/n5796 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U210  ( .ZN(\REGF/pbmemout1/n5878 ), .A(
        \pk_rread_h[20] ), .B(\pk_s8ba_h[9] ), .C(\pk_rread_h[21] ), .D(
        \pk_s7ba_h[9] ), .E(\pk_rread_h[22] ), .F(\pk_s6ba_h[9] ), .G(
        \pk_rread_h[23] ), .H(\pk_s5ba_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U591  ( .ZN(\REGF/pbmemout1/n6183 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U380  ( .ZN(\REGF/pbmemout1/n6014 ), .A(
        \REGF/RO_PCON[30] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(
        \REGF/pk_stat_h[30] ), .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U401  ( .ZN(\REGF/pbmemout1/n6031 ), .A(
        \pk_indz_h[2] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[2] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[2] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[2] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U716  ( .ZN(\REGF/pbmemout1/n6283 ), .A(
        \REGF/RO_LLPSAS[15] ), .B(\pk_rread_h[40] ), .C(1'b0), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[15] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[15] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U731  ( .ZN(\REGF/pbmemout1/n6295 ), .A(
        \pk_s4ba_h[14] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[14] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[14] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[14] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U686  ( .ZN(\REGF/pbmemout1/n6259 ), .A(
        \pk_idcy_h[16] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[16] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[16] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[16] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U237  ( .ZN(\REGF/pbmemout1/n5900 ), .A(
        \pk_sra1_h[8] ), .B(\pk_rread_h[44] ), .C(CDOUT[8]), .D(
        \pk_rread_h[45] ), .E(CDOUT[40]), .F(\pk_rread_h[46] ), .G(CDOUT[38]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U426  ( .ZN(\REGF/pbmemout1/n6051 ), .A(
        \REGF/pk_idcy_h[28] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[28] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[28] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_oai022x1 \REGF/pbmemout1/U75  ( .ZN(\pk_ada_h[31] ), .A(
        \REGF/pbmemout1/n5741 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5742 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U115  ( .Z(\pk_pdo_h[7] ), .A(
        \REGF/pbmemout1/n5773 ), .B(\REGF/pbmemout1/n5774 ), .C(
        \REGF/pbmemout1/n5775 ), .D(\REGF/pbmemout1/n5776 ) );
    snl_or04x1 \REGF/pbmemout1/U132  ( .Z(\pk_pdo_h[24] ), .A(
        \REGF/pbmemout1/n5841 ), .B(\REGF/pbmemout1/n5842 ), .C(
        \REGF/pbmemout1/n5843 ), .D(\REGF/pbmemout1/n5844 ) );
    snl_invx05 \REGF/pbmemout1/U202  ( .ZN(\REGF/pbmemout1/n5679 ), .A(
        \REGF/RO_EACC[0] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U392  ( .ZN(\REGF/pbmemout1/n6024 ), .A(
        \pk_s0ba_h[2] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[2] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[2] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[2] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U413  ( .ZN(\REGF/pbmemout1/n5864 ), .A(
        \REGF/pbmemout1/n6040 ), .B(\REGF/pbmemout1/n6039 ), .C(
        \REGF/pbmemout1/n6038 ), .D(\REGF/pbmemout1/n6037 ) );
    snl_nand04x0 \REGF/pbmemout1/U583  ( .ZN(\REGF/pbmemout1/n5830 ), .A(
        \REGF/pbmemout1/n6176 ), .B(\REGF/pbmemout1/n6175 ), .C(
        \REGF/pbmemout1/n6174 ), .D(\REGF/pbmemout1/n6173 ) );
    snl_nand04x0 \REGF/pbmemout1/U723  ( .ZN(\REGF/pbmemout1/n5806 ), .A(
        \REGF/pbmemout1/n6288 ), .B(\REGF/pbmemout1/n6287 ), .C(
        \REGF/pbmemout1/n6286 ), .D(\REGF/pbmemout1/n6285 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U694  ( .ZN(\REGF/pbmemout1/n6265 ), .A(
        \pk_s89l_h[16] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[16] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[16] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[16] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U704  ( .ZN(\REGF/pbmemout1/n6273 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_oai022x1 \REGF/pbmemout1/U90  ( .ZN(\REGF/pbmemout1/O_LDO[14] ), .A(
        \REGF/pbmemout1/n5707 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5708 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U225  ( .ZN(\REGF/pbmemout1/n5890 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[8] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[8] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U289  ( .ZN(\REGF/pbmemout1/n5941 ), .A(
        \pk_scba_h[5] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[5] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[5] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[5] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U319  ( .ZN(\REGF/pbmemout1/n5965 ), .A(
        \REGF/RO_PSTA[19] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[4] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[34]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U434  ( .ZN(\REGF/pbmemout1/n6057 ), .A(
        \pk_s89l_h[28] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[28] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[28] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[28] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U498  ( .ZN(\REGF/pbmemout1/n5845 ), .A(
        \REGF/pbmemout1/n6108 ), .B(\REGF/pbmemout1/n6107 ), .C(
        \REGF/pbmemout1/n6106 ), .D(\REGF/pbmemout1/n6105 ) );
    snl_nand04x0 \REGF/pbmemout1/U508  ( .ZN(\REGF/pbmemout1/n5843 ), .A(
        \REGF/pbmemout1/n6116 ), .B(\REGF/pbmemout1/n6115 ), .C(
        \REGF/pbmemout1/n6114 ), .D(\REGF/pbmemout1/n6113 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U350  ( .ZN(\REGF/pbmemout1/n5990 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_nand04x0 \REGF/pbmemout1/U638  ( .ZN(\REGF/pbmemout1/n5821 ), .A(
        \REGF/pbmemout1/n6220 ), .B(\REGF/pbmemout1/n6219 ), .C(
        \REGF/pbmemout1/n6218 ), .D(\REGF/pbmemout1/n6217 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U671  ( .ZN(\REGF/pbmemout1/n6247 ), .A(
        \pk_s4ba_h[17] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[17] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[17] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[17] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U541  ( .ZN(\REGF/pbmemout1/n6143 ), .A(
        \pk_indz_h[23] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[23] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[23] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[23] ), .H(\pk_rread_h[59] ) );
    snl_invx05 \REGF/pbmemout1/U147  ( .ZN(\REGF/pbmemout1/n5691 ), .A(
        \REGF/RO_ACC[6] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U377  ( .ZN(\REGF/pbmemout1/n6012 ), .A(
        \pk_sra1_h[30] ), .B(\pk_rread_h[44] ), .C(CDOUT[30]), .D(
        \pk_rread_h[45] ), .E(1'b0), .F(\pk_rread_h[46] ), .G(CDOUT[58]), .H(
        \pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U566  ( .ZN(\REGF/pbmemout1/n6163 ), .A(
        \pk_idcy_h[21] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[21] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[21] ), .F(\pk_rread_h[10] ), .G(1'b0), 
        .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U656  ( .ZN(\REGF/pbmemout1/n6235 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[18] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[18] ), .H(
        \pk_rread_h[43] ) );
    snl_nand04x0 \REGF/pbmemout1/U828  ( .ZN(\REGF/pbmemout1/n5747 ), .A(
        \REGF/pbmemout1/n6372 ), .B(\REGF/pbmemout1/n6371 ), .C(
        \REGF/pbmemout1/n6370 ), .D(\REGF/pbmemout1/n6369 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U277  ( .ZN(\REGF/pbmemout1/n5932 ), .A(
        \pk_sra1_h[6] ), .B(\pk_rread_h[44] ), .C(CDOUT[6]), .D(
        \pk_rread_h[45] ), .E(CDOUT[38]), .F(\pk_rread_h[46] ), .G(CDOUT[36]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U756  ( .ZN(\REGF/pbmemout1/n6315 ), .A(
        \REGF/RO_LLPSAS[13] ), .B(\pk_rread_h[40] ), .C(1'b0), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[13] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[13] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U814  ( .ZN(\REGF/pbmemout1/n6361 ), .A(
        \pk_s89l_h[10] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[10] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[10] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[10] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U466  ( .ZN(\REGF/pbmemout1/n6083 ), .A(
        \REGF/pk_idcy_h[26] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[26] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[26] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_invx05 \REGF/pbmemout1/U160  ( .ZN(\REGF/pbmemout1/n5738 ), .A(
        \REGF/RO_EACC[29] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U250  ( .ZN(\REGF/pbmemout1/n5910 ), .A(
        \pk_s8ba_h[7] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[7] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[7] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[7] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U441  ( .ZN(\REGF/pbmemout1/n6063 ), .A(
        \REGF/pk_indz_h[28] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[28] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[28] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[28] ), .H(\pk_rread_h[59] ) );
    snl_nand04x0 \REGF/pbmemout1/U833  ( .ZN(\REGF/pbmemout1/n5748 ), .A(
        \REGF/pbmemout1/n6376 ), .B(\REGF/pbmemout1/n6375 ), .C(
        \REGF/pbmemout1/n6374 ), .D(\REGF/pbmemout1/n6373 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U771  ( .ZN(\REGF/pbmemout1/n6327 ), .A(
        \pk_s4ba_h[12] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[12] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[12] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[12] ), .H(\pk_rread_h[27] ) );
    snl_ao222x1 \REGF/pbmemout1/U10  ( .Z(\pk_adb_h[7] ), .A(\REGF/RO_EACC[7] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[7] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[7] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U15  ( .Z(\pk_adb_h[31] ), .A(
        \REGF/RO_EACC[31] ), .B(eaccbsel), .C(\REGF/RO_SRDA[31] ), .D(
        ph_dregsl_h), .E(pk_sign_h), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U20  ( .Z(\pk_adb_h[27] ), .A(
        \REGF/RO_EACC[27] ), .B(eaccbsel), .C(\REGF/RO_SRDA[27] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[27] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U49  ( .ZN(\pk_ada_h[5] ), .A(
        \REGF/pbmemout1/n5689 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5690 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U129  ( .Z(\pk_pdo_h[21] ), .A(
        \REGF/pbmemout1/n5829 ), .B(\REGF/pbmemout1/n5830 ), .C(
        \REGF/pbmemout1/n5831 ), .D(\REGF/pbmemout1/n5832 ) );
    snl_invx05 \REGF/pbmemout1/U185  ( .ZN(\REGF/pbmemout1/n5715 ), .A(
        \REGF/RO_ACC[18] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U325  ( .ZN(\REGF/pbmemout1/n5970 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[3] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[3] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U534  ( .ZN(\REGF/pbmemout1/n6137 ), .A(
        \pk_s89l_h[23] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[23] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[23] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[23] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U292  ( .ZN(\REGF/pbmemout1/n5944 ), .A(
        \pk_s0ba_h[5] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[5] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[5] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[5] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U302  ( .ZN(\REGF/pbmemout1/n5952 ), .A(
        \pk_spr_h[5] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[5] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[5] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[5] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U483  ( .ZN(\REGF/pbmemout1/n5850 ), .A(
        \REGF/pbmemout1/n6096 ), .B(\REGF/pbmemout1/n6095 ), .C(
        \REGF/pbmemout1/n6094 ), .D(\REGF/pbmemout1/n6093 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U604  ( .ZN(\REGF/pbmemout1/n6193 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(\REGF/pk_exco_h[1] ), .D(\pk_rread_h[1] ), 
        .E(\REGF/pk_scti_h[1] ), .F(\pk_rread_h[2] ), .G(\pk_sati_h[1] ), .H(
        \pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U623  ( .ZN(\REGF/pbmemout1/n5750 ), .A(
        \REGF/pbmemout1/n6208 ), .B(\REGF/pbmemout1/n6207 ), .C(
        \REGF/pbmemout1/n6206 ), .D(\REGF/pbmemout1/n6205 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U794  ( .ZN(\REGF/pbmemout1/n6345 ), .A(
        \pk_s89l_h[11] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[11] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[11] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[11] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U513  ( .ZN(\REGF/pbmemout1/n5844 ), .A(
        \REGF/pbmemout1/n6120 ), .B(\REGF/pbmemout1/n6119 ), .C(
        \REGF/pbmemout1/n6118 ), .D(\REGF/pbmemout1/n6117 ) );
    snl_nand04x0 \REGF/pbmemout1/U738  ( .ZN(\REGF/pbmemout1/n5801 ), .A(
        \REGF/pbmemout1/n6300 ), .B(\REGF/pbmemout1/n6299 ), .C(
        \REGF/pbmemout1/n6298 ), .D(\REGF/pbmemout1/n6297 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U219  ( .ZN(\REGF/pbmemout1/n5885 ), .A(
        \pk_rread_h[48] ), .B(ph_ixco_h), .C(\pk_rread_h[49] ), .D(
        \REGF/RO_PSASL[9] ), .E(\pk_rread_h[50] ), .F(CDOUT[39]), .G(
        \pk_rread_h[51] ), .H(1'b0) );
    snl_aoi2222x0 \REGF/pbmemout1/U389  ( .ZN(\REGF/pbmemout1/n6021 ), .A(
        \pk_scba_h[2] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[2] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[2] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[2] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U408  ( .ZN(\REGF/pbmemout1/n5863 ), .A(
        \REGF/pbmemout1/n6036 ), .B(\REGF/pbmemout1/n6035 ), .C(
        \REGF/pbmemout1/n6034 ), .D(\REGF/pbmemout1/n6033 ) );
    snl_nand04x0 \REGF/pbmemout1/U598  ( .ZN(\REGF/pbmemout1/n5825 ), .A(
        \REGF/pbmemout1/n6188 ), .B(\REGF/pbmemout1/n6187 ), .C(
        \REGF/pbmemout1/n6186 ), .D(\REGF/pbmemout1/n6185 ) );
    snl_oai022x1 \REGF/pbmemout1/U69  ( .ZN(\pk_ada_h[25] ), .A(
        \REGF/pbmemout1/n5729 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5730 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U109  ( .Z(\pk_pdo_h[1] ), .A(
        \REGF/pbmemout1/n5749 ), .B(\REGF/pbmemout1/n5750 ), .C(
        \REGF/pbmemout1/n5751 ), .D(\REGF/pbmemout1/n5752 ) );
    snl_invx05 \REGF/pbmemout1/U182  ( .ZN(\REGF/pbmemout1/n5718 ), .A(
        \REGF/RO_EACC[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U295  ( .ZN(\REGF/pbmemout1/n5946 ), .A(
        \pk_s01l_h[5] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[5] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[5] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[5] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U305  ( .ZN(\REGF/pbmemout1/n5954 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[4] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[4] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U514  ( .ZN(\REGF/pbmemout1/n6121 ), .A(
        \pk_s89l_h[24] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[24] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[24] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[24] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U484  ( .ZN(\REGF/pbmemout1/n6097 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U603  ( .ZN(\REGF/pbmemout1/n5826 ), .A(
        \REGF/pbmemout1/n6192 ), .B(\REGF/pbmemout1/n6191 ), .C(
        \REGF/pbmemout1/n6190 ), .D(\REGF/pbmemout1/n6189 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U624  ( .ZN(\REGF/pbmemout1/n6209 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U793  ( .ZN(\REGF/pbmemout1/n5792 ), .A(
        \REGF/pbmemout1/n6344 ), .B(\REGF/pbmemout1/n6343 ), .C(
        \REGF/pbmemout1/n6342 ), .D(\REGF/pbmemout1/n6341 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U322  ( .ZN(\REGF/pbmemout1/n5968 ), .A(
        \pk_spr_h[4] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[4] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[4] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[4] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U533  ( .ZN(\REGF/pbmemout1/n5840 ), .A(
        \REGF/pbmemout1/n6136 ), .B(\REGF/pbmemout1/n6135 ), .C(
        \REGF/pbmemout1/n6134 ), .D(\REGF/pbmemout1/n6133 ) );
    snl_nand04x0 \REGF/pbmemout1/U688  ( .ZN(\REGF/pbmemout1/n5811 ), .A(
        \REGF/pbmemout1/n6260 ), .B(\REGF/pbmemout1/n6259 ), .C(
        \REGF/pbmemout1/n6258 ), .D(\REGF/pbmemout1/n6257 ) );
    snl_nand04x0 \REGF/pbmemout1/U718  ( .ZN(\REGF/pbmemout1/n5805 ), .A(
        \REGF/pbmemout1/n6284 ), .B(\REGF/pbmemout1/n6283 ), .C(
        \REGF/pbmemout1/n6282 ), .D(\REGF/pbmemout1/n6281 ) );
    snl_invx05 \REGF/pbmemout1/U167  ( .ZN(\REGF/pbmemout1/n5731 ), .A(
        \REGF/RO_ACC[26] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U239  ( .ZN(\REGF/pbmemout1/n5901 ), .A(
        ph_iwco_h), .B(\pk_rread_h[48] ), .C(\REGF/RO_PSASL[8] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[38]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U428  ( .ZN(\REGF/pbmemout1/n5859 ), .A(
        \REGF/pbmemout1/n6052 ), .B(\REGF/pbmemout1/n6051 ), .C(
        \REGF/pbmemout1/n6050 ), .D(\REGF/pbmemout1/n6049 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U257  ( .ZN(\REGF/pbmemout1/n5916 ), .A(
        \pk_sra1_h[7] ), .B(\pk_rread_h[44] ), .C(CDOUT[7]), .D(
        \pk_rread_h[45] ), .E(CDOUT[39]), .F(\pk_rread_h[46] ), .G(CDOUT[37]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U776  ( .ZN(\REGF/pbmemout1/n6331 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[12] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[12] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U446  ( .ZN(\REGF/pbmemout1/n6067 ), .A(
        \REGF/pk_idcy_h[27] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[27] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[27] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U834  ( .ZN(\REGF/pbmemout1/n6377 ), .A(
        \pk_s89l_h[0] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[0] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[0] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[0] ), .H(\pk_rread_h[35] ) );
    snl_ao222x1 \REGF/pbmemout1/U29  ( .Z(\pk_adb_h[19] ), .A(
        \REGF/RO_EACC[19] ), .B(eaccbsel), .C(\REGF/RO_SRDA[19] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[19] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U47  ( .ZN(\pk_ada_h[3] ), .A(
        \REGF/pbmemout1/n5685 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5686 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U55  ( .ZN(\pk_ada_h[11] ), .A(
        \REGF/pbmemout1/n5701 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5702 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U72  ( .ZN(\pk_ada_h[28] ), .A(
        \REGF/pbmemout1/n5735 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5736 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U97  ( .ZN(\REGF/pbmemout1/O_LDO[21] ), .A(
        \REGF/pbmemout1/n5721 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5722 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U140  ( .ZN(\REGF/pbmemout1/n5698 ), .A(
        \REGF/RO_EACC[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U270  ( .ZN(\REGF/pbmemout1/n5926 ), .A(
        \pk_s8ba_h[6] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[6] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[6] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[6] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U461  ( .ZN(\REGF/pbmemout1/n6079 ), .A(
        \REGF/pk_indz_h[27] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[27] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[27] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[27] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U751  ( .ZN(\REGF/pbmemout1/n6311 ), .A(
        \pk_s4ba_h[13] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[13] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[13] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[13] ), .H(\pk_rread_h[27] ) );
    snl_nand04x0 \REGF/pbmemout1/U813  ( .ZN(\REGF/pbmemout1/n5788 ), .A(
        \REGF/pbmemout1/n6360 ), .B(\REGF/pbmemout1/n6359 ), .C(
        \REGF/pbmemout1/n6358 ), .D(\REGF/pbmemout1/n6357 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U370  ( .ZN(\REGF/pbmemout1/n6006 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U651  ( .ZN(\REGF/pbmemout1/n6231 ), .A(
        \REGF/pk_s4ba_h[18] ), .B(\pk_rread_h[24] ), .C(\REGF/pk_s3ba_h[18] ), 
        .D(\pk_rread_h[25] ), .E(\REGF/pk_s2ba_h[18] ), .F(\pk_rread_h[26] ), 
        .G(\REGF/pk_s1ba_h[18] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U561  ( .ZN(\REGF/pbmemout1/n6159 ), .A(
        \pk_indz_h[22] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[22] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[22] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[22] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U222  ( .ZN(\REGF/pbmemout1/n5888 ), .A(
        \pk_rread_h[60] ), .B(\pk_spr_h[9] ), .C(\pk_rread_h[61] ), .D(
        \pk_dpr_h[9] ), .E(\pk_rread_h[62] ), .F(\REGF/RO_EACC[9] ), .G(
        \pk_rread_h[63] ), .H(\REGF/RO_ACC[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U357  ( .ZN(\REGF/pbmemout1/n5996 ), .A(
        \pk_sra1_h[31] ), .B(\pk_rread_h[44] ), .C(CDOUT[31]), .D(
        \pk_rread_h[45] ), .E(1'b0), .F(\pk_rread_h[46] ), .G(CDOUT[59]), .H(
        \pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U546  ( .ZN(\REGF/pbmemout1/n6147 ), .A(
        \pk_idcy_h[22] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[22] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[22] ), .F(\pk_rread_h[10] ), .G(1'b0), 
        .H(\pk_rread_h[11] ) );
    snl_nand04x0 \REGF/pbmemout1/U433  ( .ZN(\REGF/pbmemout1/n5860 ), .A(
        \REGF/pbmemout1/n6056 ), .B(\REGF/pbmemout1/n6055 ), .C(
        \REGF/pbmemout1/n6054 ), .D(\REGF/pbmemout1/n6053 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U676  ( .ZN(\REGF/pbmemout1/n6251 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[17] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[17] ), .H(
        \pk_rread_h[43] ) );
    snl_nand04x0 \REGF/pbmemout1/U808  ( .ZN(\REGF/pbmemout1/n5787 ), .A(
        \REGF/pbmemout1/n6356 ), .B(\REGF/pbmemout1/n6355 ), .C(
        \REGF/pbmemout1/n6354 ), .D(\REGF/pbmemout1/n6353 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U841  ( .ZN(\REGF/pbmemout1/n6383 ), .A(
        \pk_indz_h[0] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[0] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[0] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[0] ), .H(\pk_rread_h[59] ) );
    snl_or04x1 \REGF/pbmemout1/U112  ( .Z(\pk_pdo_h[4] ), .A(
        \REGF/pbmemout1/n5761 ), .B(\REGF/pbmemout1/n5762 ), .C(
        \REGF/pbmemout1/n5763 ), .D(\REGF/pbmemout1/n5764 ) );
    snl_nand04x0 \REGF/pbmemout1/U693  ( .ZN(\REGF/pbmemout1/n5812 ), .A(
        \REGF/pbmemout1/n6264 ), .B(\REGF/pbmemout1/n6263 ), .C(
        \REGF/pbmemout1/n6262 ), .D(\REGF/pbmemout1/n6261 ) );
    snl_nand04x0 \REGF/pbmemout1/U703  ( .ZN(\REGF/pbmemout1/n5810 ), .A(
        \REGF/pbmemout1/n6272 ), .B(\REGF/pbmemout1/n6271 ), .C(
        \REGF/pbmemout1/n6270 ), .D(\REGF/pbmemout1/n6269 ) );
    snl_or04x1 \REGF/pbmemout1/U135  ( .Z(\pk_pdo_h[27] ), .A(
        \REGF/pbmemout1/n5853 ), .B(\REGF/pbmemout1/n5854 ), .C(
        \REGF/pbmemout1/n5855 ), .D(\REGF/pbmemout1/n5856 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U205  ( .ZN(\REGF/pbmemout1/n5874 ), .A(
        \pk_rread_h[4] ), .B(1'b0), .C(\pk_rread_h[5] ), .D(1'b0), .E(
        \pk_rread_h[6] ), .F(\pk_saco_lh[9] ), .G(\pk_rread_h[7] ), .H(
        \pk_idcz_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U724  ( .ZN(\REGF/pbmemout1/n6289 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U395  ( .ZN(\REGF/pbmemout1/n6026 ), .A(
        \pk_s01l_h[2] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[2] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[2] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U584  ( .ZN(\REGF/pbmemout1/n6177 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U414  ( .ZN(\REGF/pbmemout1/n6041 ), .A(
        \pk_s89l_h[29] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[29] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[29] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[29] ), .H(\pk_rread_h[35] ) );
    snl_oai022x1 \REGF/pbmemout1/U60  ( .ZN(\pk_ada_h[16] ), .A(
        \REGF/pbmemout1/n5711 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5712 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_invx05 \REGF/pbmemout1/U199  ( .ZN(\REGF/pbmemout1/n5701 ), .A(
        \REGF/RO_ACC[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U339  ( .ZN(\REGF/pbmemout1/n5981 ), .A(
        \REGF/RO_PSTA[18] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[3] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[33]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U528  ( .ZN(\REGF/pbmemout1/n5839 ), .A(
        \REGF/pbmemout1/n6132 ), .B(\REGF/pbmemout1/n6131 ), .C(
        \REGF/pbmemout1/n6130 ), .D(\REGF/pbmemout1/n6129 ) );
    snl_nand04x0 \REGF/pbmemout1/U618  ( .ZN(\REGF/pbmemout1/n5749 ), .A(
        \REGF/pbmemout1/n6204 ), .B(\REGF/pbmemout1/n6203 ), .C(
        \REGF/pbmemout1/n6202 ), .D(\REGF/pbmemout1/n6201 ) );
    snl_nand04x0 \REGF/pbmemout1/U788  ( .ZN(\REGF/pbmemout1/n5791 ), .A(
        \REGF/pbmemout1/n6340 ), .B(\REGF/pbmemout1/n6339 ), .C(
        \REGF/pbmemout1/n6338 ), .D(\REGF/pbmemout1/n6337 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U230  ( .ZN(\REGF/pbmemout1/n5894 ), .A(
        \pk_s8ba_h[8] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[8] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[8] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[8] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U421  ( .ZN(\REGF/pbmemout1/n6047 ), .A(
        \REGF/pk_indz_h[29] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[29] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[29] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[29] ), .H(\pk_rread_h[59] ) );
    snl_oai022x1 \REGF/pbmemout1/U100  ( .ZN(\REGF/pbmemout1/O_LDO[24] ), .A(
        \REGF/pbmemout1/n5727 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5728 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U681  ( .ZN(\REGF/pbmemout1/n6255 ), .A(
        \pk_indz_h[17] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[17] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[17] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[17] ), .H(\pk_rread_h[59] ) );
    snl_or04x1 \REGF/pbmemout1/U127  ( .Z(\pk_pdo_h[19] ), .A(
        \REGF/pbmemout1/n5821 ), .B(\REGF/pbmemout1/n5822 ), .C(
        \REGF/pbmemout1/n5823 ), .D(\REGF/pbmemout1/n5824 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U711  ( .ZN(\REGF/pbmemout1/n6279 ), .A(
        \pk_s4ba_h[15] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[15] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[15] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[15] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U736  ( .ZN(\REGF/pbmemout1/n6299 ), .A(
        \REGF/RO_LLPSAS[14] ), .B(\pk_rread_h[40] ), .C(1'b0), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[14] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[14] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U217  ( .ZN(\REGF/pbmemout1/n5884 ), .A(
        \pk_rread_h[44] ), .B(\pk_sra1_h[9] ), .C(\pk_rread_h[45] ), .D(CDOUT
        [9]), .E(\pk_rread_h[46] ), .F(CDOUT[41]), .G(\pk_rread_h[47] ), .H(
        CDOUT[39]) );
    snl_aoi2222x0 \REGF/pbmemout1/U387  ( .ZN(\REGF/pbmemout1/n6020 ), .A(
        \pk_pcs1_h[2] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[2] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[2] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[2] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U406  ( .ZN(\REGF/pbmemout1/n6035 ), .A(
        \REGF/pk_idcy_h[29] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[29] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[29] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U596  ( .ZN(\REGF/pbmemout1/n6187 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[20] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[20] ), .H(
        \pk_rread_h[43] ) );
    snl_invx05 \REGF/pbmemout1/U149  ( .ZN(\REGF/pbmemout1/n5689 ), .A(
        \REGF/RO_ACC[5] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U279  ( .ZN(\REGF/pbmemout1/n5933 ), .A(
        \REGF/RO_EST2[6] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[6] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[36]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U758  ( .ZN(\REGF/pbmemout1/n5797 ), .A(
        \REGF/pbmemout1/n6316 ), .B(\REGF/pbmemout1/n6315 ), .C(
        \REGF/pbmemout1/n6314 ), .D(\REGF/pbmemout1/n6313 ) );
    snl_nand04x0 \REGF/pbmemout1/U468  ( .ZN(\REGF/pbmemout1/n5851 ), .A(
        \REGF/pbmemout1/n6084 ), .B(\REGF/pbmemout1/n6083 ), .C(
        \REGF/pbmemout1/n6082 ), .D(\REGF/pbmemout1/n6081 ) );
    snl_oai022x1 \REGF/pbmemout1/U85  ( .ZN(\REGF/pbmemout1/O_LDO[9] ), .A(
        \REGF/pbmemout1/n5697 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5698 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U362  ( .ZN(\REGF/pbmemout1/n6000 ), .A(
        \pk_spr_h[31] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[31] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[31] ), .F(\pk_rread_h[62] ), .G(
        pk_sign_h), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U573  ( .ZN(\REGF/pbmemout1/n5832 ), .A(
        \REGF/pbmemout1/n6168 ), .B(\REGF/pbmemout1/n6167 ), .C(
        \REGF/pbmemout1/n6166 ), .D(\REGF/pbmemout1/n6165 ) );
    snl_nand04x0 \REGF/pbmemout1/U643  ( .ZN(\REGF/pbmemout1/n5822 ), .A(
        \REGF/pbmemout1/n6224 ), .B(\REGF/pbmemout1/n6223 ), .C(
        \REGF/pbmemout1/n6222 ), .D(\REGF/pbmemout1/n6221 ) );
    snl_invx05 \REGF/pbmemout1/U175  ( .ZN(\REGF/pbmemout1/n5723 ), .A(
        \REGF/RO_ACC[22] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U345  ( .ZN(\REGF/pbmemout1/n5986 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_hh[31] ), .F(\pk_rread_h[6] ), .G(\REGF/pk_idcz_h[31] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U379  ( .ZN(\REGF/pbmemout1/n6013 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[58]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U554  ( .ZN(\REGF/pbmemout1/n6153 ), .A(
        \pk_s89l_h[22] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[22] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[22] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[22] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U568  ( .ZN(\REGF/pbmemout1/n5831 ), .A(
        \REGF/pbmemout1/n6164 ), .B(\REGF/pbmemout1/n6163 ), .C(
        \REGF/pbmemout1/n6162 ), .D(\REGF/pbmemout1/n6161 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U664  ( .ZN(\REGF/pbmemout1/n6241 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U658  ( .ZN(\REGF/pbmemout1/n5817 ), .A(
        \REGF/pbmemout1/n6236 ), .B(\REGF/pbmemout1/n6235 ), .C(
        \REGF/pbmemout1/n6234 ), .D(\REGF/pbmemout1/n6233 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U764  ( .ZN(\REGF/pbmemout1/n6321 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_ao222x1 \REGF/pbmemout1/U17  ( .Z(\pk_adb_h[2] ), .A(\REGF/RO_EACC[2] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[2] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[2] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U22  ( .Z(\pk_adb_h[25] ), .A(
        \REGF/RO_EACC[25] ), .B(eaccbsel), .C(\REGF/RO_SRDA[25] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[25] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U32  ( .Z(\pk_adb_h[16] ), .A(
        \REGF/RO_EACC[16] ), .B(eaccbsel), .C(\REGF/RO_SRDA[16] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[16] ), .F(accbsel) );
    snl_aoi2222x0 \REGF/pbmemout1/U245  ( .ZN(\REGF/pbmemout1/n5906 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[7] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[7] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U454  ( .ZN(\REGF/pbmemout1/n6073 ), .A(
        \pk_s89l_h[27] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[27] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[27] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[27] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U826  ( .ZN(\REGF/pbmemout1/n6371 ), .A(
        \pk_idcy_h[0] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[0] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[0] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[0] ), .H(\pk_rread_h[11] ) );
    snl_ao222x1 \REGF/pbmemout1/U39  ( .Z(\pk_adb_h[0] ), .A(\REGF/RO_EACC[0] 
        ), .B(eaccbsel), .C(pk_rgbit_h), .D(ph_dregsl_h), .E(\REGF/RO_ACC[0] ), 
        .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U57  ( .ZN(\pk_ada_h[13] ), .A(
        \REGF/pbmemout1/n5705 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5706 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U137  ( .Z(\pk_pdo_h[29] ), .A(
        \REGF/pbmemout1/n5861 ), .B(\REGF/pbmemout1/n5862 ), .C(
        \REGF/pbmemout1/n5863 ), .D(\REGF/pbmemout1/n5864 ) );
    snl_invx05 \REGF/pbmemout1/U152  ( .ZN(\REGF/pbmemout1/n5686 ), .A(
        \REGF/RO_EACC[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U262  ( .ZN(\REGF/pbmemout1/n5920 ), .A(
        \pk_spr_h[7] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[7] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[7] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[7] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U801  ( .ZN(\REGF/pbmemout1/n6351 ), .A(
        \pk_indz_h[11] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[11] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[11] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[11] ), .H(\pk_rread_h[59] ) );
    snl_nand04x0 \REGF/pbmemout1/U473  ( .ZN(\REGF/pbmemout1/n5852 ), .A(
        \REGF/pbmemout1/n6088 ), .B(\REGF/pbmemout1/n6087 ), .C(
        \REGF/pbmemout1/n6086 ), .D(\REGF/pbmemout1/n6085 ) );
    snl_invx05 \REGF/pbmemout1/U190  ( .ZN(\REGF/pbmemout1/n5710 ), .A(
        \REGF/RO_EACC[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U287  ( .ZN(\REGF/pbmemout1/n5940 ), .A(
        \pk_pcs1_h[5] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[5] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[5] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[5] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U317  ( .ZN(\REGF/pbmemout1/n5964 ), .A(
        \pk_sra1_h[4] ), .B(\pk_rread_h[44] ), .C(CDOUT[4]), .D(
        \pk_rread_h[45] ), .E(CDOUT[36]), .F(\pk_rread_h[46] ), .G(CDOUT[34]), 
        .H(\pk_rread_h[47] ) );
    snl_nand04x0 \REGF/pbmemout1/U743  ( .ZN(\REGF/pbmemout1/n5802 ), .A(
        \REGF/pbmemout1/n6304 ), .B(\REGF/pbmemout1/n6303 ), .C(
        \REGF/pbmemout1/n6302 ), .D(\REGF/pbmemout1/n6301 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U496  ( .ZN(\REGF/pbmemout1/n6107 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[25] ), .F(\pk_rread_h[42] ), .G(1'b0), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U506  ( .ZN(\REGF/pbmemout1/n6115 ), .A(
        \REGF/pk_idcy_h[24] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[24] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[24] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U611  ( .ZN(\REGF/pbmemout1/n6199 ), .A(
        \pk_s4ba_h[1] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[1] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[1] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[1] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U636  ( .ZN(\REGF/pbmemout1/n6219 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[19] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[19] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U330  ( .ZN(\REGF/pbmemout1/n5974 ), .A(
        \pk_s8ba_h[3] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[3] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[3] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[3] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U521  ( .ZN(\REGF/pbmemout1/n6127 ), .A(
        \REGF/pk_indz_h[24] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[24] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[24] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[24] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U781  ( .ZN(\REGF/pbmemout1/n6335 ), .A(
        \pk_indz_h[12] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[12] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[12] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[12] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U726  ( .ZN(\REGF/pbmemout1/n6291 ), .A(
        \pk_idcy_h[14] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[14] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[14] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[14] ), .H(\pk_rread_h[11] ) );
    snl_oai022x1 \REGF/pbmemout1/U70  ( .ZN(\pk_ada_h[26] ), .A(
        \REGF/pbmemout1/n5731 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5732 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U207  ( .ZN(\REGF/pbmemout1/n5876 ), .A(
        \pk_rread_h[12] ), .B(\pk_pcs1_h[9] ), .C(\pk_rread_h[13] ), .D(
        \pk_sfba_h[9] ), .E(\pk_rread_h[14] ), .F(\pk_seba_h[9] ), .G(
        \pk_rread_h[15] ), .H(\pk_sdba_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U397  ( .ZN(\REGF/pbmemout1/n6028 ), .A(
        \pk_sra1_h[2] ), .B(\pk_rread_h[44] ), .C(CDOUT[2]), .D(
        \pk_rread_h[45] ), .E(CDOUT[34]), .F(\pk_rread_h[46] ), .G(CDOUT[32]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U586  ( .ZN(\REGF/pbmemout1/n6179 ), .A(
        \pk_idcy_h[20] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[20] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[20] ), .F(\pk_rread_h[10] ), .G(1'b0), 
        .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U416  ( .ZN(\REGF/pbmemout1/n6043 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[29] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[29] ), .H(
        \pk_rread_h[43] ) );
    snl_or04x1 \REGF/pbmemout1/U110  ( .Z(\pk_pdo_h[2] ), .A(
        \REGF/pbmemout1/n5753 ), .B(\REGF/pbmemout1/n5754 ), .C(
        \REGF/pbmemout1/n5755 ), .D(\REGF/pbmemout1/n5756 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U220  ( .ZN(\REGF/pbmemout1/n5886 ), .A(
        \pk_rread_h[52] ), .B(\REGF/RO_PCON[9] ), .C(\pk_rread_h[53] ), .D(
        \REGF/RO_PPCN[9] ), .E(\pk_rread_h[54] ), .F(\pk_pc_h[9] ), .G(
        \pk_rread_h[55] ), .H(1'b0) );
    snl_aoi2222x0 \REGF/pbmemout1/U431  ( .ZN(\REGF/pbmemout1/n6055 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_nand04x0 \REGF/pbmemout1/U843  ( .ZN(\REGF/pbmemout1/n5746 ), .A(
        \REGF/pbmemout1/n6384 ), .B(\REGF/pbmemout1/n6383 ), .C(
        \REGF/pbmemout1/n6382 ), .D(\REGF/pbmemout1/n6381 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U691  ( .ZN(\REGF/pbmemout1/n6263 ), .A(
        \pk_s4ba_h[16] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[16] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[16] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[16] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U701  ( .ZN(\REGF/pbmemout1/n6271 ), .A(
        \pk_indz_h[16] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[16] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[16] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[16] ), .H(\pk_rread_h[59] ) );
    snl_invx05 \REGF/pbmemout1/U159  ( .ZN(\REGF/pbmemout1/n5683 ), .A(
        \REGF/RO_ACC[2] ) );
    snl_nand04x0 \REGF/pbmemout1/U748  ( .ZN(\REGF/pbmemout1/n5799 ), .A(
        \REGF/pbmemout1/n6308 ), .B(\REGF/pbmemout1/n6307 ), .C(
        \REGF/pbmemout1/n6306 ), .D(\REGF/pbmemout1/n6305 ) );
    snl_oai022x1 \REGF/pbmemout1/U95  ( .ZN(\REGF/pbmemout1/O_LDO[19] ), .A(
        \REGF/pbmemout1/n5717 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5718 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U269  ( .ZN(\REGF/pbmemout1/n5925 ), .A(
        \pk_scba_h[6] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[6] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[6] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[6] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U478  ( .ZN(\REGF/pbmemout1/n5849 ), .A(
        \REGF/pbmemout1/n6092 ), .B(\REGF/pbmemout1/n6091 ), .C(
        \REGF/pbmemout1/n6090 ), .D(\REGF/pbmemout1/n6089 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U355  ( .ZN(\REGF/pbmemout1/n5994 ), .A(
        \pk_s01l_h[31] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[31] ), .F(\pk_rread_h[38] ), .G(1'b0), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U544  ( .ZN(\REGF/pbmemout1/n6145 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U272  ( .ZN(\REGF/pbmemout1/n5928 ), .A(
        \pk_s0ba_h[6] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[6] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[6] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[6] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U369  ( .ZN(\REGF/pbmemout1/n6005 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U372  ( .ZN(\REGF/pbmemout1/n6008 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[30] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[30] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[30] ), .H(
        \pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U653  ( .ZN(\REGF/pbmemout1/n5820 ), .A(
        \REGF/pbmemout1/n6232 ), .B(\REGF/pbmemout1/n6231 ), .C(
        \REGF/pbmemout1/n6230 ), .D(\REGF/pbmemout1/n6229 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U674  ( .ZN(\REGF/pbmemout1/n6249 ), .A(
        \pk_s89l_h[17] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[17] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[17] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[17] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U563  ( .ZN(\REGF/pbmemout1/n5834 ), .A(
        \REGF/pbmemout1/n6160 ), .B(\REGF/pbmemout1/n6159 ), .C(
        \REGF/pbmemout1/n6158 ), .D(\REGF/pbmemout1/n6157 ) );
    snl_nand04x0 \REGF/pbmemout1/U463  ( .ZN(\REGF/pbmemout1/n5854 ), .A(
        \REGF/pbmemout1/n6080 ), .B(\REGF/pbmemout1/n6079 ), .C(
        \REGF/pbmemout1/n6078 ), .D(\REGF/pbmemout1/n6077 ) );
    snl_nand04x0 \REGF/pbmemout1/U578  ( .ZN(\REGF/pbmemout1/n5829 ), .A(
        \REGF/pbmemout1/n6172 ), .B(\REGF/pbmemout1/n6171 ), .C(
        \REGF/pbmemout1/n6170 ), .D(\REGF/pbmemout1/n6169 ) );
    snl_nand04x0 \REGF/pbmemout1/U648  ( .ZN(\REGF/pbmemout1/n5819 ), .A(
        \REGF/pbmemout1/n6228 ), .B(\REGF/pbmemout1/n6227 ), .C(
        \REGF/pbmemout1/n6226 ), .D(\REGF/pbmemout1/n6225 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U811  ( .ZN(\REGF/pbmemout1/n6359 ), .A(
        \pk_s4ba_h[10] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[10] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[10] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[10] ), .H(\pk_rread_h[27] ) );
    snl_ao222x1 \REGF/pbmemout1/U30  ( .Z(\pk_adb_h[18] ), .A(
        \REGF/RO_EACC[18] ), .B(eaccbsel), .C(\REGF/RO_SRDA[18] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[18] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U79  ( .ZN(\REGF/pbmemout1/O_LDO[3] ), .A(
        \REGF/pbmemout1/n5685 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5686 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U119  ( .Z(\pk_pdo_h[11] ), .A(
        \REGF/pbmemout1/n5789 ), .B(\REGF/pbmemout1/n5790 ), .C(
        \REGF/pbmemout1/n5791 ), .D(\REGF/pbmemout1/n5792 ) );
    snl_invx05 \REGF/pbmemout1/U142  ( .ZN(\REGF/pbmemout1/n5696 ), .A(
        \REGF/RO_EACC[8] ) );
    snl_nand04x0 \REGF/pbmemout1/U753  ( .ZN(\REGF/pbmemout1/n5800 ), .A(
        \REGF/pbmemout1/n6312 ), .B(\REGF/pbmemout1/n6311 ), .C(
        \REGF/pbmemout1/n6310 ), .D(\REGF/pbmemout1/n6309 ) );
    snl_invx05 \REGF/pbmemout1/U165  ( .ZN(\REGF/pbmemout1/n5733 ), .A(
        \REGF/RO_ACC[27] ) );
    snl_invx05 \REGF/pbmemout1/U180  ( .ZN(\REGF/pbmemout1/n5682 ), .A(
        \REGF/RO_EACC[1] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U255  ( .ZN(\REGF/pbmemout1/n5914 ), .A(
        \pk_s01l_h[7] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[7] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[7] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[7] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U774  ( .ZN(\REGF/pbmemout1/n6329 ), .A(
        \pk_s89l_h[12] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[12] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[12] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[12] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U836  ( .ZN(\REGF/pbmemout1/n6379 ), .A(
        \REGF/RO_LLPSAS[0] ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[0] ), .D(
        \pk_rread_h[41] ), .E(pk_rgbit_h), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[0] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U444  ( .ZN(\REGF/pbmemout1/n6065 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U601  ( .ZN(\REGF/pbmemout1/n6191 ), .A(
        \pk_indz_h[20] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[20] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[20] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[20] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U791  ( .ZN(\REGF/pbmemout1/n6343 ), .A(
        \pk_s4ba_h[11] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[11] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[11] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[11] ), .H(\pk_rread_h[27] ) );
    snl_invx05 \REGF/pbmemout1/U192  ( .ZN(\REGF/pbmemout1/n5708 ), .A(
        \REGF/RO_EACC[14] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U297  ( .ZN(\REGF/pbmemout1/n5948 ), .A(
        \pk_sra1_h[5] ), .B(\pk_rread_h[44] ), .C(CDOUT[5]), .D(
        \pk_rread_h[45] ), .E(CDOUT[37]), .F(\pk_rread_h[46] ), .G(CDOUT[35]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U320  ( .ZN(\REGF/pbmemout1/n5966 ), .A(
        \REGF/RO_PCON[4] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[4] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[4] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U531  ( .ZN(\REGF/pbmemout1/n6135 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U307  ( .ZN(\REGF/pbmemout1/n5956 ), .A(
        \pk_pcs1_h[4] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[4] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[4] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[4] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U516  ( .ZN(\REGF/pbmemout1/n6123 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[24] ), .F(\pk_rread_h[42] ), .G(1'b0), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U486  ( .ZN(\REGF/pbmemout1/n6099 ), .A(
        \REGF/pk_idcy_h[25] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[25] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[25] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_nand04x0 \REGF/pbmemout1/U613  ( .ZN(\REGF/pbmemout1/n5752 ), .A(
        \REGF/pbmemout1/n6200 ), .B(\REGF/pbmemout1/n6199 ), .C(
        \REGF/pbmemout1/n6198 ), .D(\REGF/pbmemout1/n6197 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U626  ( .ZN(\REGF/pbmemout1/n6211 ), .A(
        \pk_idcy_h[19] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[19] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[19] ), .F(\pk_rread_h[10] ), .G(1'b0), 
        .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U285  ( .ZN(\REGF/pbmemout1/n5938 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[5] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[5] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U315  ( .ZN(\REGF/pbmemout1/n5962 ), .A(
        \pk_s01l_h[4] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[4] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[4] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[4] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U332  ( .ZN(\REGF/pbmemout1/n5976 ), .A(
        \pk_s0ba_h[3] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[3] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[3] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[3] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U523  ( .ZN(\REGF/pbmemout1/n5842 ), .A(
        \REGF/pbmemout1/n6128 ), .B(\REGF/pbmemout1/n6127 ), .C(
        \REGF/pbmemout1/n6126 ), .D(\REGF/pbmemout1/n6125 ) );
    snl_nand04x0 \REGF/pbmemout1/U783  ( .ZN(\REGF/pbmemout1/n5794 ), .A(
        \REGF/pbmemout1/n6336 ), .B(\REGF/pbmemout1/n6335 ), .C(
        \REGF/pbmemout1/n6334 ), .D(\REGF/pbmemout1/n6333 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U494  ( .ZN(\REGF/pbmemout1/n6105 ), .A(
        \pk_s89l_h[25] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[25] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[25] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[25] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U504  ( .ZN(\REGF/pbmemout1/n6113 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U634  ( .ZN(\REGF/pbmemout1/n6217 ), .A(
        \pk_s89l_h[19] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[19] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[19] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[19] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U698  ( .ZN(\REGF/pbmemout1/n5809 ), .A(
        \REGF/pbmemout1/n6268 ), .B(\REGF/pbmemout1/n6267 ), .C(
        \REGF/pbmemout1/n6266 ), .D(\REGF/pbmemout1/n6265 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U229  ( .ZN(\REGF/pbmemout1/n5893 ), .A(
        \pk_scba_h[8] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[8] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[8] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[8] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U708  ( .ZN(\REGF/pbmemout1/n5807 ), .A(
        \REGF/pbmemout1/n6276 ), .B(\REGF/pbmemout1/n6275 ), .C(
        \REGF/pbmemout1/n6274 ), .D(\REGF/pbmemout1/n6273 ) );
    snl_nand04x0 \REGF/pbmemout1/U438  ( .ZN(\REGF/pbmemout1/n5857 ), .A(
        \REGF/pbmemout1/n6060 ), .B(\REGF/pbmemout1/n6059 ), .C(
        \REGF/pbmemout1/n6058 ), .D(\REGF/pbmemout1/n6057 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U260  ( .ZN(\REGF/pbmemout1/n5918 ), .A(
        \REGF/RO_PCON[7] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[7] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[7] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U471  ( .ZN(\REGF/pbmemout1/n6087 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_nand04x0 \REGF/pbmemout1/U803  ( .ZN(\REGF/pbmemout1/n5790 ), .A(
        \REGF/pbmemout1/n6352 ), .B(\REGF/pbmemout1/n6351 ), .C(
        \REGF/pbmemout1/n6350 ), .D(\REGF/pbmemout1/n6349 ) );
    snl_invx05 \REGF/pbmemout1/U150  ( .ZN(\REGF/pbmemout1/n5688 ), .A(
        \REGF/RO_EACC[4] ) );
    snl_invx05 \REGF/pbmemout1/U177  ( .ZN(\REGF/pbmemout1/n5721 ), .A(
        \REGF/RO_ACC[21] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U741  ( .ZN(\REGF/pbmemout1/n6303 ), .A(
        \pk_indz_h[14] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[14] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[14] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[14] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U766  ( .ZN(\REGF/pbmemout1/n6323 ), .A(
        \pk_idcy_h[12] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[12] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[12] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[12] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U247  ( .ZN(\REGF/pbmemout1/n5908 ), .A(
        \pk_pcs1_h[7] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[7] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[7] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[7] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U456  ( .ZN(\REGF/pbmemout1/n6075 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[27] ), .F(\pk_rread_h[42] ), .G(1'b0), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U824  ( .ZN(\REGF/pbmemout1/n6369 ), .A(
        \REGF/RO_ERFA[0] ), .B(\pk_rread_h[0] ), .C(\REGF/pk_exco_h[0] ), .D(
        \pk_rread_h[1] ), .E(\REGF/pk_scti_h[0] ), .F(\pk_rread_h[2] ), .G(
        \pk_sati_h[0] ), .H(\pk_rread_h[3] ) );
    snl_invx1 \REGF/pbmemout1/U42  ( .ZN(\REGF/pbmemout1/n5744 ), .A(
        po_reacl_h) );
    snl_oai022x1 \REGF/pbmemout1/U45  ( .ZN(\pk_ada_h[1] ), .A(
        \REGF/pbmemout1/n5681 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5682 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U87  ( .ZN(\REGF/pbmemout1/O_LDO[11] ), .A(
        \REGF/pbmemout1/n5701 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5702 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U347  ( .ZN(\REGF/pbmemout1/n5988 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U556  ( .ZN(\REGF/pbmemout1/n6155 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[22] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[22] ), .H(
        \pk_rread_h[43] ) );
    snl_or04x1 \REGF/pbmemout1/U125  ( .Z(\pk_pdo_h[17] ), .A(
        \REGF/pbmemout1/n5813 ), .B(\REGF/pbmemout1/n5814 ), .C(
        \REGF/pbmemout1/n5815 ), .D(\REGF/pbmemout1/n5816 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U360  ( .ZN(\REGF/pbmemout1/n5998 ), .A(
        pk_pcon31_h), .B(\pk_rread_h[52] ), .C(1'b0), .D(\pk_rread_h[53] ), 
        .E(1'b0), .F(\pk_rread_h[54] ), .G(\REGF/pk_stat_h[31] ), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U571  ( .ZN(\REGF/pbmemout1/n6167 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U641  ( .ZN(\REGF/pbmemout1/n6223 ), .A(
        \pk_indz_h[19] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[19] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[19] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[19] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U666  ( .ZN(\REGF/pbmemout1/n6243 ), .A(
        \pk_idcy_h[17] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[17] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[17] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[17] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U734  ( .ZN(\REGF/pbmemout1/n6297 ), .A(
        \pk_s89l_h[14] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[14] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[14] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[14] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U818  ( .ZN(\REGF/pbmemout1/n5785 ), .A(
        \REGF/pbmemout1/n6364 ), .B(\REGF/pbmemout1/n6363 ), .C(
        \REGF/pbmemout1/n6362 ), .D(\REGF/pbmemout1/n6361 ) );
    snl_oai022x1 \REGF/pbmemout1/U62  ( .ZN(\pk_ada_h[18] ), .A(
        \REGF/pbmemout1/n5715 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5716 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U215  ( .ZN(\REGF/pbmemout1/n5882 ), .A(
        \pk_rread_h[36] ), .B(\pk_s01l_h[9] ), .C(\pk_rread_h[37] ), .D(
        \pk_stdat[9] ), .E(\pk_rread_h[38] ), .F(\pk_trba_h[9] ), .G(
        \pk_rread_h[39] ), .H(\REGF/RO_ERRA[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U385  ( .ZN(\REGF/pbmemout1/n6018 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[2] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[2] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U404  ( .ZN(\REGF/pbmemout1/n6033 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U594  ( .ZN(\REGF/pbmemout1/n6185 ), .A(
        \pk_s89l_h[20] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[20] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[20] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[20] ), .H(\pk_rread_h[35] ) );
    snl_oai022x1 \REGF/pbmemout1/U65  ( .ZN(\pk_ada_h[21] ), .A(
        \REGF/pbmemout1/n5721 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5722 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U102  ( .ZN(\REGF/pbmemout1/O_LDO[26] ), .A(
        \REGF/pbmemout1/n5731 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5732 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U232  ( .ZN(\REGF/pbmemout1/n5896 ), .A(
        \pk_s0ba_h[8] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[8] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[8] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[8] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U423  ( .ZN(\REGF/pbmemout1/n5862 ), .A(
        \REGF/pbmemout1/n6048 ), .B(\REGF/pbmemout1/n6047 ), .C(
        \REGF/pbmemout1/n6046 ), .D(\REGF/pbmemout1/n6045 ) );
    snl_nand04x0 \REGF/pbmemout1/U683  ( .ZN(\REGF/pbmemout1/n5814 ), .A(
        \REGF/pbmemout1/n6256 ), .B(\REGF/pbmemout1/n6255 ), .C(
        \REGF/pbmemout1/n6254 ), .D(\REGF/pbmemout1/n6253 ) );
    snl_oai022x1 \REGF/pbmemout1/U105  ( .ZN(\REGF/pbmemout1/O_LDO[29] ), .A(
        \REGF/pbmemout1/n5737 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5738 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U189  ( .ZN(\REGF/pbmemout1/n5711 ), .A(
        \REGF/RO_ACC[16] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U329  ( .ZN(\REGF/pbmemout1/n5973 ), .A(
        \pk_scba_h[3] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[3] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[3] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[3] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U538  ( .ZN(\REGF/pbmemout1/n5837 ), .A(
        \REGF/pbmemout1/n6140 ), .B(\REGF/pbmemout1/n6139 ), .C(
        \REGF/pbmemout1/n6138 ), .D(\REGF/pbmemout1/n6137 ) );
    snl_nand04x0 \REGF/pbmemout1/U713  ( .ZN(\REGF/pbmemout1/n5808 ), .A(
        \REGF/pbmemout1/n6280 ), .B(\REGF/pbmemout1/n6279 ), .C(
        \REGF/pbmemout1/n6278 ), .D(\REGF/pbmemout1/n6277 ) );
    snl_nand04x0 \REGF/pbmemout1/U608  ( .ZN(\REGF/pbmemout1/n5751 ), .A(
        \REGF/pbmemout1/n6196 ), .B(\REGF/pbmemout1/n6195 ), .C(
        \REGF/pbmemout1/n6194 ), .D(\REGF/pbmemout1/n6193 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U714  ( .ZN(\REGF/pbmemout1/n6281 ), .A(
        \pk_s89l_h[15] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[15] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[15] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[15] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U798  ( .ZN(\REGF/pbmemout1/n5789 ), .A(
        \REGF/pbmemout1/n6348 ), .B(\REGF/pbmemout1/n6347 ), .C(
        \REGF/pbmemout1/n6346 ), .D(\REGF/pbmemout1/n6345 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U235  ( .ZN(\REGF/pbmemout1/n5898 ), .A(
        \pk_s01l_h[8] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[8] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[8] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[8] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U424  ( .ZN(\REGF/pbmemout1/n6049 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U684  ( .ZN(\REGF/pbmemout1/n6257 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U212  ( .ZN(\REGF/pbmemout1/n5880 ), .A(
        \pk_rread_h[28] ), .B(\pk_s0ba_h[9] ), .C(\pk_rread_h[29] ), .D(
        \pk_sefl_h[9] ), .E(\pk_rread_h[30] ), .F(\pk_scdl_h[9] ), .G(
        \pk_rread_h[31] ), .H(\pk_sabl_h[9] ) );
    snl_nand04x0 \REGF/pbmemout1/U593  ( .ZN(\REGF/pbmemout1/n5828 ), .A(
        \REGF/pbmemout1/n6184 ), .B(\REGF/pbmemout1/n6183 ), .C(
        \REGF/pbmemout1/n6182 ), .D(\REGF/pbmemout1/n6181 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U382  ( .ZN(\REGF/pbmemout1/n6016 ), .A(
        \pk_spr_h[30] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[30] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[30] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[30] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U403  ( .ZN(\REGF/pbmemout1/n5754 ), .A(
        \REGF/pbmemout1/n6032 ), .B(\REGF/pbmemout1/n6031 ), .C(
        \REGF/pbmemout1/n6030 ), .D(\REGF/pbmemout1/n6029 ) );
    snl_oai022x1 \REGF/pbmemout1/U80  ( .ZN(\REGF/pbmemout1/O_LDO[4] ), .A(
        \REGF/pbmemout1/n5687 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5688 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U122  ( .Z(\pk_pdo_h[14] ), .A(
        \REGF/pbmemout1/n5801 ), .B(\REGF/pbmemout1/n5802 ), .C(
        \REGF/pbmemout1/n5803 ), .D(\REGF/pbmemout1/n5804 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U299  ( .ZN(\REGF/pbmemout1/n5949 ), .A(
        \REGF/RO_EST2[5] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[5] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[35]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U518  ( .ZN(\REGF/pbmemout1/n5841 ), .A(
        \REGF/pbmemout1/n6124 ), .B(\REGF/pbmemout1/n6123 ), .C(
        \REGF/pbmemout1/n6122 ), .D(\REGF/pbmemout1/n6121 ) );
    snl_nand04x0 \REGF/pbmemout1/U733  ( .ZN(\REGF/pbmemout1/n5804 ), .A(
        \REGF/pbmemout1/n6296 ), .B(\REGF/pbmemout1/n6295 ), .C(
        \REGF/pbmemout1/n6294 ), .D(\REGF/pbmemout1/n6293 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U309  ( .ZN(\REGF/pbmemout1/n5957 ), .A(
        \pk_scba_h[4] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[4] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[4] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[4] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U488  ( .ZN(\REGF/pbmemout1/n5847 ), .A(
        \REGF/pbmemout1/n6100 ), .B(\REGF/pbmemout1/n6099 ), .C(
        \REGF/pbmemout1/n6098 ), .D(\REGF/pbmemout1/n6097 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U367  ( .ZN(\REGF/pbmemout1/n6004 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_nand04x0 \REGF/pbmemout1/U628  ( .ZN(\REGF/pbmemout1/n5823 ), .A(
        \REGF/pbmemout1/n6212 ), .B(\REGF/pbmemout1/n6211 ), .C(
        \REGF/pbmemout1/n6210 ), .D(\REGF/pbmemout1/n6209 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U576  ( .ZN(\REGF/pbmemout1/n6171 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[21] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[21] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U646  ( .ZN(\REGF/pbmemout1/n6227 ), .A(
        \pk_idcy_h[18] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[18] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[18] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[18] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U661  ( .ZN(\REGF/pbmemout1/n6239 ), .A(
        \pk_indz_h[18] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[18] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[18] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[18] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U340  ( .ZN(\REGF/pbmemout1/n5982 ), .A(
        \REGF/RO_PCON[3] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[3] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[3] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U551  ( .ZN(\REGF/pbmemout1/n6151 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_nand04x0 \REGF/pbmemout1/U838  ( .ZN(\REGF/pbmemout1/n5745 ), .A(
        \REGF/pbmemout1/n6380 ), .B(\REGF/pbmemout1/n6379 ), .C(
        \REGF/pbmemout1/n6378 ), .D(\REGF/pbmemout1/n6377 ) );
    snl_ao222x1 \REGF/pbmemout1/U11  ( .Z(\pk_adb_h[6] ), .A(\REGF/RO_EACC[6] 
        ), .B(eaccbsel), .C(\REGF/RO_SRDA[6] ), .D(ph_dregsl_h), .E(
        \REGF/RO_ACC[6] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U19  ( .Z(\pk_adb_h[28] ), .A(
        \REGF/RO_EACC[28] ), .B(eaccbsel), .C(\REGF/RO_SRDA[28] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[28] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U25  ( .Z(\pk_adb_h[22] ), .A(
        \REGF/RO_EACC[22] ), .B(eaccbsel), .C(\REGF/RO_SRDA[22] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[22] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U37  ( .Z(\pk_adb_h[11] ), .A(
        \REGF/RO_EACC[11] ), .B(eaccbsel), .C(\REGF/RO_SRDA[11] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[11] ), .F(accbsel) );
    snl_invx05 \REGF/pbmemout1/U157  ( .ZN(\REGF/pbmemout1/n5739 ), .A(
        \REGF/RO_ACC[30] ) );
    snl_invx05 \REGF/pbmemout1/U170  ( .ZN(\REGF/pbmemout1/n5728 ), .A(
        \REGF/RO_EACC[24] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U240  ( .ZN(\REGF/pbmemout1/n5902 ), .A(
        \REGF/RO_PCON[8] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[8] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[8] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_nand04x0 \REGF/pbmemout1/U823  ( .ZN(\REGF/pbmemout1/n5786 ), .A(
        \REGF/pbmemout1/n6368 ), .B(\REGF/pbmemout1/n6367 ), .C(
        \REGF/pbmemout1/n6366 ), .D(\REGF/pbmemout1/n6365 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U451  ( .ZN(\REGF/pbmemout1/n6071 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U746  ( .ZN(\REGF/pbmemout1/n6307 ), .A(
        \pk_idcy_h[13] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[13] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[13] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[13] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U761  ( .ZN(\REGF/pbmemout1/n6319 ), .A(
        \pk_indz_h[13] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[13] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[13] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[13] ), .H(\pk_rread_h[59] ) );
    snl_oai022x1 \REGF/pbmemout1/U59  ( .ZN(\pk_ada_h[15] ), .A(
        \REGF/pbmemout1/n5709 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5710 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U139  ( .Z(\pk_pdo_h[31] ), .A(
        \REGF/pbmemout1/n5869 ), .B(\REGF/pbmemout1/n5870 ), .C(
        \REGF/pbmemout1/n5871 ), .D(\REGF/pbmemout1/n5872 ) );
    snl_invx05 \REGF/pbmemout1/U195  ( .ZN(\REGF/pbmemout1/n5705 ), .A(
        \REGF/RO_ACC[13] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U267  ( .ZN(\REGF/pbmemout1/n5924 ), .A(
        \pk_pcs1_h[6] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[6] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[6] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[6] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U476  ( .ZN(\REGF/pbmemout1/n6091 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[26] ), .F(\pk_rread_h[42] ), .G(1'b0), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U804  ( .ZN(\REGF/pbmemout1/n6353 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U282  ( .ZN(\REGF/pbmemout1/n5936 ), .A(
        \pk_spr_h[6] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[6] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[6] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[6] ), .H(\pk_rread_h[63] ) );
    snl_nand04x0 \REGF/pbmemout1/U503  ( .ZN(\REGF/pbmemout1/n5846 ), .A(
        \REGF/pbmemout1/n6112 ), .B(\REGF/pbmemout1/n6111 ), .C(
        \REGF/pbmemout1/n6110 ), .D(\REGF/pbmemout1/n6109 ) );
    snl_nand04x0 \REGF/pbmemout1/U633  ( .ZN(\REGF/pbmemout1/n5824 ), .A(
        \REGF/pbmemout1/n6216 ), .B(\REGF/pbmemout1/n6215 ), .C(
        \REGF/pbmemout1/n6214 ), .D(\REGF/pbmemout1/n6213 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U312  ( .ZN(\REGF/pbmemout1/n5960 ), .A(
        \pk_s0ba_h[4] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[4] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[4] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[4] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U493  ( .ZN(\REGF/pbmemout1/n5848 ), .A(
        \REGF/pbmemout1/n6104 ), .B(\REGF/pbmemout1/n6103 ), .C(
        \REGF/pbmemout1/n6102 ), .D(\REGF/pbmemout1/n6101 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U335  ( .ZN(\REGF/pbmemout1/n5978 ), .A(
        \pk_s01l_h[3] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[3] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[3] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U524  ( .ZN(\REGF/pbmemout1/n6129 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U784  ( .ZN(\REGF/pbmemout1/n6337 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U614  ( .ZN(\REGF/pbmemout1/n6201 ), .A(
        \pk_s89l_h[1] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[1] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[1] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[1] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U728  ( .ZN(\REGF/pbmemout1/n5803 ), .A(
        \REGF/pbmemout1/n6292 ), .B(\REGF/pbmemout1/n6291 ), .C(
        \REGF/pbmemout1/n6290 ), .D(\REGF/pbmemout1/n6289 ) );
    snl_oai022x1 \REGF/pbmemout1/U89  ( .ZN(\REGF/pbmemout1/O_LDO[13] ), .A(
        \REGF/pbmemout1/n5705 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5706 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_invx05 \REGF/pbmemout1/U187  ( .ZN(\REGF/pbmemout1/n5713 ), .A(
        \REGF/RO_ACC[17] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U209  ( .ZN(\REGF/pbmemout1/n5877 ), .A(
        \pk_rread_h[16] ), .B(\pk_scba_h[9] ), .C(\pk_rread_h[17] ), .D(
        \pk_sbba_h[9] ), .E(\pk_rread_h[18] ), .F(\pk_saba_h[9] ), .G(
        \pk_rread_h[19] ), .H(\pk_s9ba_h[9] ) );
    snl_nand04x0 \REGF/pbmemout1/U588  ( .ZN(\REGF/pbmemout1/n5827 ), .A(
        \REGF/pbmemout1/n6180 ), .B(\REGF/pbmemout1/n6179 ), .C(
        \REGF/pbmemout1/n6178 ), .D(\REGF/pbmemout1/n6177 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U290  ( .ZN(\REGF/pbmemout1/n5942 ), .A(
        \pk_s8ba_h[5] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[5] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[5] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[5] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U300  ( .ZN(\REGF/pbmemout1/n5950 ), .A(
        \REGF/RO_PCON[5] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[5] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[5] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U399  ( .ZN(\REGF/pbmemout1/n6029 ), .A(
        \REGF/RO_EST2[2] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[2] ), .D(
        \pk_rread_h[49] ), .E(CDOUT[32]), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U418  ( .ZN(\REGF/pbmemout1/n5861 ), .A(
        \REGF/pbmemout1/n6044 ), .B(\REGF/pbmemout1/n6043 ), .C(
        \REGF/pbmemout1/n6042 ), .D(\REGF/pbmemout1/n6041 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U481  ( .ZN(\REGF/pbmemout1/n6095 ), .A(
        \REGF/pk_indz_h[26] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[26] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[26] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[26] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U621  ( .ZN(\REGF/pbmemout1/n6207 ), .A(
        \pk_indz_h[1] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[1] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[1] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[1] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U511  ( .ZN(\REGF/pbmemout1/n6119 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U327  ( .ZN(\REGF/pbmemout1/n5972 ), .A(
        \pk_pcs1_h[3] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[3] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[3] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[3] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U536  ( .ZN(\REGF/pbmemout1/n6139 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[23] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[23] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U349  ( .ZN(\REGF/pbmemout1/n5989 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U606  ( .ZN(\REGF/pbmemout1/n6195 ), .A(
        \pk_idcy_h[1] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[1] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[1] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[1] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U796  ( .ZN(\REGF/pbmemout1/n6347 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[11] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[11] ), .H(
        \pk_rread_h[43] ) );
    snl_nand04x0 \REGF/pbmemout1/U558  ( .ZN(\REGF/pbmemout1/n5833 ), .A(
        \REGF/pbmemout1/n6156 ), .B(\REGF/pbmemout1/n6155 ), .C(
        \REGF/pbmemout1/n6154 ), .D(\REGF/pbmemout1/n6153 ) );
    snl_invx05 \REGF/pbmemout1/U145  ( .ZN(\REGF/pbmemout1/n5693 ), .A(
        \REGF/RO_ACC[7] ) );
    snl_invx05 \REGF/pbmemout1/U162  ( .ZN(\REGF/pbmemout1/n5736 ), .A(
        \REGF/RO_EACC[28] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U252  ( .ZN(\REGF/pbmemout1/n5912 ), .A(
        \pk_s0ba_h[7] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[7] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[7] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[7] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U443  ( .ZN(\REGF/pbmemout1/n5858 ), .A(
        \REGF/pbmemout1/n6064 ), .B(\REGF/pbmemout1/n6063 ), .C(
        \REGF/pbmemout1/n6062 ), .D(\REGF/pbmemout1/n6061 ) );
    snl_nand04x0 \REGF/pbmemout1/U668  ( .ZN(\REGF/pbmemout1/n5815 ), .A(
        \REGF/pbmemout1/n6244 ), .B(\REGF/pbmemout1/n6243 ), .C(
        \REGF/pbmemout1/n6242 ), .D(\REGF/pbmemout1/n6241 ) );
    snl_nand04x0 \REGF/pbmemout1/U773  ( .ZN(\REGF/pbmemout1/n5796 ), .A(
        \REGF/pbmemout1/n6328 ), .B(\REGF/pbmemout1/n6327 ), .C(
        \REGF/pbmemout1/n6326 ), .D(\REGF/pbmemout1/n6325 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U831  ( .ZN(\REGF/pbmemout1/n6375 ), .A(
        \pk_s4ba_h[0] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[0] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[0] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[0] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U754  ( .ZN(\REGF/pbmemout1/n6313 ), .A(
        \pk_s89l_h[13] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[13] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[13] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[13] ), .H(\pk_rread_h[35] ) );
    snl_invx05 \REGF/pbmemout1/U179  ( .ZN(\REGF/pbmemout1/n5719 ), .A(
        \REGF/RO_ACC[20] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U275  ( .ZN(\REGF/pbmemout1/n5930 ), .A(
        \pk_s01l_h[6] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[6] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[6] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[6] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U464  ( .ZN(\REGF/pbmemout1/n6081 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U768  ( .ZN(\REGF/pbmemout1/n5795 ), .A(
        \REGF/pbmemout1/n6324 ), .B(\REGF/pbmemout1/n6323 ), .C(
        \REGF/pbmemout1/n6322 ), .D(\REGF/pbmemout1/n6321 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U816  ( .ZN(\REGF/pbmemout1/n6363 ), .A(
        \REGF/RO_LLPSAS[10] ), .B(\pk_rread_h[40] ), .C(1'b0), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[10] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[10] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U249  ( .ZN(\REGF/pbmemout1/n5909 ), .A(
        \pk_scba_h[7] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[7] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[7] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[7] ), .H(\pk_rread_h[19] ) );
    snl_nand04x0 \REGF/pbmemout1/U458  ( .ZN(\REGF/pbmemout1/n5853 ), .A(
        \REGF/pbmemout1/n6076 ), .B(\REGF/pbmemout1/n6075 ), .C(
        \REGF/pbmemout1/n6074 ), .D(\REGF/pbmemout1/n6073 ) );
    snl_oai022x1 \REGF/pbmemout1/U50  ( .ZN(\pk_ada_h[6] ), .A(
        \REGF/pbmemout1/n5691 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5692 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U77  ( .ZN(\REGF/pbmemout1/O_LDO[1] ), .A(
        \REGF/pbmemout1/n5681 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5682 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_oai022x1 \REGF/pbmemout1/U92  ( .ZN(\REGF/pbmemout1/O_LDO[16] ), .A(
        \REGF/pbmemout1/n5711 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5712 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U375  ( .ZN(\REGF/pbmemout1/n6010 ), .A(
        \pk_s01l_h[30] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[30] ), .F(\pk_rread_h[38] ), .G(1'b0), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U564  ( .ZN(\REGF/pbmemout1/n6161 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(1'b0), .F(
        \pk_rread_h[2] ), .G(1'b0), .H(\pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U654  ( .ZN(\REGF/pbmemout1/n6233 ), .A(
        \pk_s89l_h[18] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[18] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[18] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[18] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U673  ( .ZN(\REGF/pbmemout1/n5816 ), .A(
        \REGF/pbmemout1/n6248 ), .B(\REGF/pbmemout1/n6247 ), .C(
        \REGF/pbmemout1/n6246 ), .D(\REGF/pbmemout1/n6245 ) );
    snl_or04x1 \REGF/pbmemout1/U117  ( .Z(\pk_pdo_h[9] ), .A(
        \REGF/pbmemout1/n5781 ), .B(\REGF/pbmemout1/n5782 ), .C(
        \REGF/pbmemout1/n5783 ), .D(\REGF/pbmemout1/n5784 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U352  ( .ZN(\REGF/pbmemout1/n5992 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[31] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[31] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[31] ), .H(
        \pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U543  ( .ZN(\REGF/pbmemout1/n5838 ), .A(
        \REGF/pbmemout1/n6144 ), .B(\REGF/pbmemout1/n6143 ), .C(
        \REGF/pbmemout1/n6142 ), .D(\REGF/pbmemout1/n6141 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U227  ( .ZN(\REGF/pbmemout1/n5892 ), .A(
        \pk_pcs1_h[8] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[8] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[8] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[8] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U696  ( .ZN(\REGF/pbmemout1/n6267 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[16] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[16] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U706  ( .ZN(\REGF/pbmemout1/n6275 ), .A(
        \pk_idcy_h[15] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[15] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[15] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[15] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U436  ( .ZN(\REGF/pbmemout1/n6059 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(1'b0), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[28] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[28] ), .H(
        \pk_rread_h[43] ) );
    snl_invx05 \REGF/pbmemout1/U200  ( .ZN(\REGF/pbmemout1/n5700 ), .A(
        \REGF/RO_EACC[10] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U390  ( .ZN(\REGF/pbmemout1/n6022 ), .A(
        \pk_s8ba_h[2] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[2] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[2] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[2] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U411  ( .ZN(\REGF/pbmemout1/n6039 ), .A(1'b0
        ), .B(\pk_rread_h[24] ), .C(1'b0), .D(\pk_rread_h[25] ), .E(1'b0), .F(
        \pk_rread_h[26] ), .G(1'b0), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U581  ( .ZN(\REGF/pbmemout1/n6175 ), .A(
        \pk_indz_h[21] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[21] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[21] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[21] ), .H(\pk_rread_h[59] ) );
    snl_oai022x1 \REGF/pbmemout1/U58  ( .ZN(\pk_ada_h[14] ), .A(
        \REGF/pbmemout1/n5707 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5708 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_or04x1 \REGF/pbmemout1/U130  ( .Z(\pk_pdo_h[22] ), .A(
        \REGF/pbmemout1/n5833 ), .B(\REGF/pbmemout1/n5834 ), .C(
        \REGF/pbmemout1/n5835 ), .D(\REGF/pbmemout1/n5836 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U721  ( .ZN(\REGF/pbmemout1/n6287 ), .A(
        \pk_indz_h[15] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[15] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[15] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[15] ), .H(\pk_rread_h[59] ) );
    snl_or04x1 \REGF/pbmemout1/U138  ( .Z(\pk_pdo_h[30] ), .A(
        \REGF/pbmemout1/n5865 ), .B(\REGF/pbmemout1/n5866 ), .C(
        \REGF/pbmemout1/n5867 ), .D(\REGF/pbmemout1/n5868 ) );
    snl_invx05 \REGF/pbmemout1/U194  ( .ZN(\REGF/pbmemout1/n5706 ), .A(
        \REGF/RO_EACC[13] ) );
    snl_nand04x0 \REGF/pbmemout1/U283  ( .ZN(\REGF/pbmemout1/n5770 ), .A(
        \REGF/pbmemout1/n5936 ), .B(\REGF/pbmemout1/n5935 ), .C(
        \REGF/pbmemout1/n5934 ), .D(\REGF/pbmemout1/n5933 ) );
    snl_nand04x0 \REGF/pbmemout1/U313  ( .ZN(\REGF/pbmemout1/n5764 ), .A(
        \REGF/pbmemout1/n5960 ), .B(\REGF/pbmemout1/n5959 ), .C(
        \REGF/pbmemout1/n5958 ), .D(\REGF/pbmemout1/n5957 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U632  ( .ZN(\REGF/pbmemout1/n6216 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[19] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[19] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[19] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U492  ( .ZN(\REGF/pbmemout1/n6104 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[25] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[25] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[25] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U334  ( .ZN(\REGF/pbmemout1/n5977 ), .A(
        \pk_s89l_h[3] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[3] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[3] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[3] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U502  ( .ZN(\REGF/pbmemout1/n6112 ), .A(1'b0
        ), .B(\pk_rread_h[60] ), .C(1'b0), .D(\pk_rread_h[61] ), .E(
        \REGF/RO_EACC[25] ), .F(\pk_rread_h[62] ), .G(\REGF/RO_ACC[25] ), .H(
        \pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U525  ( .ZN(\REGF/pbmemout1/n6130 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[23] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[23] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U615  ( .ZN(\REGF/pbmemout1/n6202 ), .A(
        \pk_s01l_h[1] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[1] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[1] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U729  ( .ZN(\REGF/pbmemout1/n6293 ), .A(
        \pk_scba_h[14] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[14] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[14] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[14] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U785  ( .ZN(\REGF/pbmemout1/n6338 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[11] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[11] ), .H(
        \pk_rread_h[7] ) );
    snl_nand04x0 \REGF/pbmemout1/U208  ( .ZN(\REGF/pbmemout1/n5783 ), .A(
        \REGF/pbmemout1/n5876 ), .B(\REGF/pbmemout1/n5875 ), .C(
        \REGF/pbmemout1/n5874 ), .D(\REGF/pbmemout1/n5873 ) );
    snl_nand04x0 \REGF/pbmemout1/U398  ( .ZN(\REGF/pbmemout1/n5753 ), .A(
        \REGF/pbmemout1/n6028 ), .B(\REGF/pbmemout1/n6027 ), .C(
        \REGF/pbmemout1/n6026 ), .D(\REGF/pbmemout1/n6025 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U419  ( .ZN(\REGF/pbmemout1/n6045 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[57]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U589  ( .ZN(\REGF/pbmemout1/n6181 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U241  ( .ZN(\REGF/pbmemout1/n5903 ), .A(
        \pk_indz_h[8] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[8] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[8] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[8] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U450  ( .ZN(\REGF/pbmemout1/n6070 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U822  ( .ZN(\REGF/pbmemout1/n6368 ), .A(
        \pk_spr_h[10] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[10] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[10] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[10] ), .H(\pk_rread_h[63] ) );
    snl_ao222x1 \REGF/pbmemout1/U16  ( .Z(\pk_adb_h[30] ), .A(
        \REGF/RO_EACC[30] ), .B(eaccbsel), .C(\REGF/RO_SRDA[30] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[30] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U18  ( .Z(\pk_adb_h[29] ), .A(
        \REGF/RO_EACC[29] ), .B(eaccbsel), .C(\REGF/RO_SRDA[29] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[29] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U36  ( .Z(\pk_adb_h[12] ), .A(
        \REGF/RO_EACC[12] ), .B(eaccbsel), .C(\REGF/RO_SRDA[12] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[12] ), .F(accbsel) );
    snl_invx05 \REGF/pbmemout1/U156  ( .ZN(\REGF/pbmemout1/n5740 ), .A(
        \REGF/RO_EACC[30] ) );
    snl_invx05 \REGF/pbmemout1/U171  ( .ZN(\REGF/pbmemout1/n5727 ), .A(
        \REGF/RO_ACC[24] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U760  ( .ZN(\REGF/pbmemout1/n6318 ), .A(
        \REGF/RO_PCON[13] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[13] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[13] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U266  ( .ZN(\REGF/pbmemout1/n5923 ), .A(
        \pk_idcy_h[6] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[6] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[6] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[6] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U747  ( .ZN(\REGF/pbmemout1/n6308 ), .A(
        \pk_pcs1_h[13] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[13] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[13] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[13] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U805  ( .ZN(\REGF/pbmemout1/n6354 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[10] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[10] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U477  ( .ZN(\REGF/pbmemout1/n6092 ), .A(1'b0
        ), .B(\pk_rread_h[44] ), .C(CDOUT[26]), .D(\pk_rread_h[45] ), .E(CDOUT
        [58]), .F(\pk_rread_h[46] ), .G(\pk_stat_h[0] ), .H(\pk_rread_h[47] )
         );
    snl_invx2 \REGF/pbmemout1/U43  ( .ZN(\REGF/pbmemout1/n5678 ), .A(accasel)
         );
    snl_oai022x1 \REGF/pbmemout1/U64  ( .ZN(\pk_ada_h[20] ), .A(
        \REGF/pbmemout1/n5719 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5720 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U81  ( .ZN(\REGF/pbmemout1/O_LDO[5] ), .A(
        \REGF/pbmemout1/n5689 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5690 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U341  ( .ZN(\REGF/pbmemout1/n5983 ), .A(
        \pk_indz_h[3] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[3] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[3] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[3] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U366  ( .ZN(\REGF/pbmemout1/n6003 ), .A(
        \REGF/pk_idcy_h[30] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[30] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[30] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U577  ( .ZN(\REGF/pbmemout1/n6172 ), .A(
        \pk_sra1_h[21] ), .B(\pk_rread_h[44] ), .C(CDOUT[21]), .D(
        \pk_rread_h[45] ), .E(CDOUT[53]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[21] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U647  ( .ZN(\REGF/pbmemout1/n6228 ), .A(
        \pk_pcs1_h[18] ), .B(\pk_rread_h[12] ), .C(\REGF/pk_sfba_h[18] ), .D(
        \pk_rread_h[13] ), .E(\REGF/pk_seba_h[18] ), .F(\pk_rread_h[14] ), .G(
        \REGF/pk_sdba_h[18] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U660  ( .ZN(\REGF/pbmemout1/n6238 ), .A(
        \REGF/RO_PCON[18] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[18] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[18] ), .F(\pk_rread_h[54] ), .G(
        \pk_stat_h[18] ), .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U550  ( .ZN(\REGF/pbmemout1/n6150 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_oai022x1 \REGF/pbmemout1/U104  ( .ZN(\REGF/pbmemout1/O_LDO[28] ), .A(
        \REGF/pbmemout1/n5735 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5736 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U685  ( .ZN(\REGF/pbmemout1/n6258 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[16] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[16] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U839  ( .ZN(\REGF/pbmemout1/n6381 ), .A(
        \REGF/RO_EST2[0] ), .B(\pk_rread_h[48] ), .C(\REGF/RO_EST1[0] ), .D(
        \pk_rread_h[49] ), .E(1'b0), .F(\pk_rread_h[50] ), .G(pk_pexe01_h), 
        .H(\pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U715  ( .ZN(\REGF/pbmemout1/n6282 ), .A(
        \pk_s01l_h[15] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[15] ), .F(\pk_rread_h[38] ), .G(\REGF/RO_ERRA[15] ), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U234  ( .ZN(\REGF/pbmemout1/n5897 ), .A(
        \pk_s89l_h[8] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[8] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[8] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[8] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U425  ( .ZN(\REGF/pbmemout1/n6050 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_hh[28] ), .F(\pk_rread_h[6] ), .G(\REGF/pk_idcz_h[28] ), .H(
        \pk_rread_h[7] ) );
    snl_oai022x1 \REGF/pbmemout1/U51  ( .ZN(\pk_ada_h[7] ), .A(
        \REGF/pbmemout1/n5693 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5694 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U76  ( .ZN(\REGF/pbmemout1/O_LDO[0] ), .A(
        \REGF/pbmemout1/n5677 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5679 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U116  ( .Z(\pk_pdo_h[8] ), .A(
        \REGF/pbmemout1/n5777 ), .B(\REGF/pbmemout1/n5778 ), .C(
        \REGF/pbmemout1/n5779 ), .D(\REGF/pbmemout1/n5780 ) );
    snl_or04x1 \REGF/pbmemout1/U123  ( .Z(\pk_pdo_h[15] ), .A(
        \REGF/pbmemout1/n5805 ), .B(\REGF/pbmemout1/n5806 ), .C(
        \REGF/pbmemout1/n5807 ), .D(\REGF/pbmemout1/n5808 ) );
    snl_nand04x0 \REGF/pbmemout1/U213  ( .ZN(\REGF/pbmemout1/n5784 ), .A(
        \REGF/pbmemout1/n5880 ), .B(\REGF/pbmemout1/n5879 ), .C(
        \REGF/pbmemout1/n5878 ), .D(\REGF/pbmemout1/n5877 ) );
    snl_nand04x0 \REGF/pbmemout1/U383  ( .ZN(\REGF/pbmemout1/n5866 ), .A(
        \REGF/pbmemout1/n6016 ), .B(\REGF/pbmemout1/n6015 ), .C(
        \REGF/pbmemout1/n6014 ), .D(\REGF/pbmemout1/n6013 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U402  ( .ZN(\REGF/pbmemout1/n6032 ), .A(
        \pk_spr_h[2] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[2] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[2] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[2] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U592  ( .ZN(\REGF/pbmemout1/n6184 ), .A(1'b0
        ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[20] ), .D(\pk_rread_h[29] ), 
        .E(\pk_scdl_h[20] ), .F(\pk_rread_h[30] ), .G(\pk_sabl_h[20] ), .H(
        \pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U732  ( .ZN(\REGF/pbmemout1/n6296 ), .A(
        \pk_s0ba_h[14] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[14] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[14] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[14] ), .H(\pk_rread_h[31] ) );
    snl_nand04x0 \REGF/pbmemout1/U298  ( .ZN(\REGF/pbmemout1/n5765 ), .A(
        \REGF/pbmemout1/n5948 ), .B(\REGF/pbmemout1/n5947 ), .C(
        \REGF/pbmemout1/n5946 ), .D(\REGF/pbmemout1/n5945 ) );
    snl_nand04x0 \REGF/pbmemout1/U308  ( .ZN(\REGF/pbmemout1/n5763 ), .A(
        \REGF/pbmemout1/n5956 ), .B(\REGF/pbmemout1/n5955 ), .C(
        \REGF/pbmemout1/n5954 ), .D(\REGF/pbmemout1/n5953 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U489  ( .ZN(\REGF/pbmemout1/n6101 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U519  ( .ZN(\REGF/pbmemout1/n6125 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/pk_stat_h[16] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U629  ( .ZN(\REGF/pbmemout1/n6213 ), .A(1'b0
        ), .B(\pk_rread_h[16] ), .C(1'b0), .D(\pk_rread_h[17] ), .E(1'b0), .F(
        \pk_rread_h[18] ), .G(1'b0), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U697  ( .ZN(\REGF/pbmemout1/n6268 ), .A(
        \pk_sra1_h[16] ), .B(\pk_rread_h[44] ), .C(CDOUT[16]), .D(
        \pk_rread_h[45] ), .E(CDOUT[48]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[16] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U707  ( .ZN(\REGF/pbmemout1/n6276 ), .A(
        \pk_pcs1_h[15] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[15] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[15] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[15] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U226  ( .ZN(\REGF/pbmemout1/n5891 ), .A(
        \pk_idcy_h[8] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[8] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[8] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[8] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U437  ( .ZN(\REGF/pbmemout1/n6060 ), .A(
        \pk_sra1_h[28] ), .B(\pk_rread_h[44] ), .C(CDOUT[28]), .D(
        \pk_rread_h[45] ), .E(1'b0), .F(\pk_rread_h[46] ), .G(CDOUT[56]), .H(
        \pk_rread_h[47] ) );
    snl_or04x1 \REGF/pbmemout1/U131  ( .Z(\pk_pdo_h[23] ), .A(
        \REGF/pbmemout1/n5837 ), .B(\REGF/pbmemout1/n5838 ), .C(
        \REGF/pbmemout1/n5839 ), .D(\REGF/pbmemout1/n5840 ) );
    snl_invx05 \REGF/pbmemout1/U201  ( .ZN(\REGF/pbmemout1/n5699 ), .A(
        \REGF/RO_ACC[10] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U391  ( .ZN(\REGF/pbmemout1/n6023 ), .A(
        \pk_s4ba_h[2] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[2] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[2] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[2] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U580  ( .ZN(\REGF/pbmemout1/n6174 ), .A(
        \REGF/RO_PCON[21] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U410  ( .ZN(\REGF/pbmemout1/n6038 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_invx05 \REGF/pbmemout1/U178  ( .ZN(\REGF/pbmemout1/n5720 ), .A(
        \REGF/RO_EACC[20] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U720  ( .ZN(\REGF/pbmemout1/n6286 ), .A(
        \REGF/RO_PCON[15] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[15] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[15] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U769  ( .ZN(\REGF/pbmemout1/n6325 ), .A(
        \pk_scba_h[12] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[12] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[12] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[12] ), .H(\pk_rread_h[19] ) );
    snl_ao222x1 \REGF/pbmemout1/U23  ( .Z(\pk_adb_h[24] ), .A(
        \REGF/RO_EACC[24] ), .B(eaccbsel), .C(\REGF/RO_SRDA[24] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[24] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U24  ( .Z(\pk_adb_h[23] ), .A(
        \REGF/RO_EACC[23] ), .B(eaccbsel), .C(\REGF/RO_SRDA[23] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[23] ), .F(accbsel) );
    snl_oai022x1 \REGF/pbmemout1/U88  ( .ZN(\REGF/pbmemout1/O_LDO[12] ), .A(
        \REGF/pbmemout1/n5703 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5704 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_oai022x1 \REGF/pbmemout1/U93  ( .ZN(\REGF/pbmemout1/O_LDO[17] ), .A(
        \REGF/pbmemout1/n5713 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5714 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_nand04x0 \REGF/pbmemout1/U248  ( .ZN(\REGF/pbmemout1/n5775 ), .A(
        \REGF/pbmemout1/n5908 ), .B(\REGF/pbmemout1/n5907 ), .C(
        \REGF/pbmemout1/n5906 ), .D(\REGF/pbmemout1/n5905 ) );
    snl_nand04x0 \REGF/pbmemout1/U353  ( .ZN(\REGF/pbmemout1/n5872 ), .A(
        \REGF/pbmemout1/n5992 ), .B(\REGF/pbmemout1/n5991 ), .C(
        \REGF/pbmemout1/n5990 ), .D(\REGF/pbmemout1/n5989 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U374  ( .ZN(\REGF/pbmemout1/n6009 ), .A(
        \pk_s89l_h[30] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[30] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[30] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[30] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U459  ( .ZN(\REGF/pbmemout1/n6077 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[55]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U542  ( .ZN(\REGF/pbmemout1/n6144 ), .A(
        \pk_spr_h[23] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[23] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[23] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[23] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U565  ( .ZN(\REGF/pbmemout1/n6162 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[21] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[21] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U655  ( .ZN(\REGF/pbmemout1/n6234 ), .A(
        \pk_s01l_h[18] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[14] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[18] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[18] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U672  ( .ZN(\REGF/pbmemout1/n6248 ), .A(
        \pk_s0ba_h[17] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[17] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[17] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[17] ), .H(\pk_rread_h[31] ) );
    snl_invx05 \REGF/pbmemout1/U144  ( .ZN(\REGF/pbmemout1/n5694 ), .A(
        \REGF/RO_EACC[7] ) );
    snl_invx05 \REGF/pbmemout1/U163  ( .ZN(\REGF/pbmemout1/n5735 ), .A(
        \REGF/RO_ACC[28] ) );
    snl_nand04x0 \REGF/pbmemout1/U253  ( .ZN(\REGF/pbmemout1/n5776 ), .A(
        \REGF/pbmemout1/n5912 ), .B(\REGF/pbmemout1/n5911 ), .C(
        \REGF/pbmemout1/n5910 ), .D(\REGF/pbmemout1/n5909 ) );
    snl_nand04x0 \REGF/pbmemout1/U348  ( .ZN(\REGF/pbmemout1/n5871 ), .A(
        \REGF/pbmemout1/n5988 ), .B(\REGF/pbmemout1/n5987 ), .C(
        \REGF/pbmemout1/n5986 ), .D(\REGF/pbmemout1/n5985 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U559  ( .ZN(\REGF/pbmemout1/n6157 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[22] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U669  ( .ZN(\REGF/pbmemout1/n6245 ), .A(
        \pk_scba_h[17] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[17] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[17] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[17] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U442  ( .ZN(\REGF/pbmemout1/n6064 ), .A(
        \pk_spr_h[28] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[28] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[28] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[28] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U830  ( .ZN(\REGF/pbmemout1/n6374 ), .A(
        \pk_s8ba_h[0] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[0] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[0] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[0] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U755  ( .ZN(\REGF/pbmemout1/n6314 ), .A(
        \pk_s01l_h[13] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[13] ), .F(\pk_rread_h[38] ), .G(\REGF/RO_ERRA[13] ), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U772  ( .ZN(\REGF/pbmemout1/n6328 ), .A(
        \pk_s0ba_h[12] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[12] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[12] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[12] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U274  ( .ZN(\REGF/pbmemout1/n5929 ), .A(
        \pk_s89l_h[6] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[6] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[6] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[6] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U465  ( .ZN(\REGF/pbmemout1/n6082 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(1'b0), .F(
        \pk_rread_h[6] ), .G(\REGF/pk_idcz_h[26] ), .H(\pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U817  ( .ZN(\REGF/pbmemout1/n6364 ), .A(
        \pk_sra1_h[10] ), .B(\pk_rread_h[44] ), .C(CDOUT[10]), .D(
        \pk_rread_h[45] ), .E(CDOUT[42]), .F(\pk_rread_h[46] ), .G(CDOUT[40]), 
        .H(\pk_rread_h[47] ) );
    snl_invx05 \REGF/pbmemout1/U181  ( .ZN(\REGF/pbmemout1/n5681 ), .A(
        \REGF/RO_ACC[1] ) );
    snl_invx05 \REGF/pbmemout1/U186  ( .ZN(\REGF/pbmemout1/n5714 ), .A(
        \REGF/RO_EACC[17] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U291  ( .ZN(\REGF/pbmemout1/n5943 ), .A(
        \pk_s4ba_h[5] ), .B(\pk_rread_h[24] ), .C(\pk_s3ba_h[5] ), .D(
        \pk_rread_h[25] ), .E(\pk_s2ba_h[5] ), .F(\pk_rread_h[26] ), .G(
        \pk_s1ba_h[5] ), .H(\pk_rread_h[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U620  ( .ZN(\REGF/pbmemout1/n6206 ), .A(
        \REGF/RO_PCON[1] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[1] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[1] ), .F(\pk_rread_h[54] ), .G(
        \pk_stat_h[1] ), .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U301  ( .ZN(\REGF/pbmemout1/n5951 ), .A(
        \pk_indz_h[5] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[5] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[5] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[5] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U510  ( .ZN(\REGF/pbmemout1/n6118 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U326  ( .ZN(\REGF/pbmemout1/n5971 ), .A(
        \pk_idcy_h[3] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[3] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[3] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[3] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U480  ( .ZN(\REGF/pbmemout1/n6094 ), .A(
        \REGF/RO_PCON[26] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U537  ( .ZN(\REGF/pbmemout1/n6140 ), .A(
        \pk_sra1_h[23] ), .B(\pk_rread_h[44] ), .C(CDOUT[23]), .D(
        \pk_rread_h[45] ), .E(CDOUT[55]), .F(\pk_rread_h[46] ), .G(
        \pk_stat_h[18] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U607  ( .ZN(\REGF/pbmemout1/n6196 ), .A(
        \pk_pcs1_h[1] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[1] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[1] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[1] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U797  ( .ZN(\REGF/pbmemout1/n6348 ), .A(
        \pk_sra1_h[11] ), .B(\pk_rread_h[44] ), .C(CDOUT[11]), .D(
        \pk_rread_h[45] ), .E(CDOUT[43]), .F(\pk_rread_h[46] ), .G(CDOUT[41]), 
        .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U296  ( .ZN(\REGF/pbmemout1/n5947 ), .A(
        \REGF/RO_LLPSAS[5] ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[5] ), .D(
        \pk_rread_h[41] ), .E(\REGF/RO_SRDA[5] ), .F(\pk_rread_h[42] ), .G(
        \pk_sra2_h[5] ), .H(\pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U306  ( .ZN(\REGF/pbmemout1/n5955 ), .A(
        \pk_idcy_h[4] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[4] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[4] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[4] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U321  ( .ZN(\REGF/pbmemout1/n5967 ), .A(
        \pk_indz_h[4] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[4] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[4] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[4] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U530  ( .ZN(\REGF/pbmemout1/n6134 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U600  ( .ZN(\REGF/pbmemout1/n6190 ), .A(
        \REGF/RO_PCON[20] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U790  ( .ZN(\REGF/pbmemout1/n6342 ), .A(
        \pk_s8ba_h[11] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[11] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[11] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[11] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U487  ( .ZN(\REGF/pbmemout1/n6100 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U517  ( .ZN(\REGF/pbmemout1/n6124 ), .A(1'b0
        ), .B(\pk_rread_h[44] ), .C(CDOUT[24]), .D(\pk_rread_h[45] ), .E(CDOUT
        [56]), .F(\pk_rread_h[46] ), .G(\REGF/pk_stat_h[16] ), .H(
        \pk_rread_h[47] ) );
    snl_nand04x0 \REGF/pbmemout1/U368  ( .ZN(\REGF/pbmemout1/n5867 ), .A(
        \REGF/pbmemout1/n6004 ), .B(\REGF/pbmemout1/n6003 ), .C(
        \REGF/pbmemout1/n6002 ), .D(\REGF/pbmemout1/n6001 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U579  ( .ZN(\REGF/pbmemout1/n6173 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[21] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U627  ( .ZN(\REGF/pbmemout1/n6212 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U649  ( .ZN(\REGF/pbmemout1/n6229 ), .A(
        \REGF/pk_scba_h[18] ), .B(\pk_rread_h[16] ), .C(\REGF/pk_sbba_h[18] ), 
        .D(\pk_rread_h[17] ), .E(\REGF/pk_saba_h[18] ), .F(\pk_rread_h[18] ), 
        .G(\REGF/pk_s9ba_h[18] ), .H(\pk_rread_h[19] ) );
    snl_ao222x1 \REGF/pbmemout1/U31  ( .Z(\pk_adb_h[17] ), .A(
        \REGF/RO_EACC[17] ), .B(eaccbsel), .C(\REGF/RO_SRDA[17] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[17] ), .F(accbsel) );
    snl_ao222x1 \REGF/pbmemout1/U38  ( .Z(\pk_adb_h[10] ), .A(
        \REGF/RO_EACC[10] ), .B(eaccbsel), .C(\REGF/RO_SRDA[10] ), .D(
        ph_dregsl_h), .E(\REGF/RO_ACC[10] ), .F(accbsel) );
    snl_invx05 \REGF/pbmemout1/U143  ( .ZN(\REGF/pbmemout1/n5695 ), .A(
        \REGF/RO_ACC[8] ) );
    snl_nand04x0 \REGF/pbmemout1/U273  ( .ZN(\REGF/pbmemout1/n5772 ), .A(
        \REGF/pbmemout1/n5928 ), .B(\REGF/pbmemout1/n5927 ), .C(
        \REGF/pbmemout1/n5926 ), .D(\REGF/pbmemout1/n5925 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U810  ( .ZN(\REGF/pbmemout1/n6358 ), .A(
        \pk_s8ba_h[10] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[10] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[10] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[10] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U462  ( .ZN(\REGF/pbmemout1/n6080 ), .A(1'b0
        ), .B(\pk_rread_h[60] ), .C(1'b0), .D(\pk_rread_h[61] ), .E(
        \REGF/RO_EACC[27] ), .F(\pk_rread_h[62] ), .G(\REGF/RO_ACC[27] ), .H(
        \pk_rread_h[63] ) );
    snl_invx05 \REGF/pbmemout1/U158  ( .ZN(\REGF/pbmemout1/n5684 ), .A(
        \REGF/RO_EACC[2] ) );
    snl_invx05 \REGF/pbmemout1/U164  ( .ZN(\REGF/pbmemout1/n5734 ), .A(
        \REGF/RO_EACC[27] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U752  ( .ZN(\REGF/pbmemout1/n6312 ), .A(
        \pk_s0ba_h[13] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[13] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[13] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[13] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U775  ( .ZN(\REGF/pbmemout1/n6330 ), .A(
        \pk_s01l_h[12] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[12] ), .F(\pk_rread_h[38] ), .G(\REGF/RO_ERRA[12] ), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U254  ( .ZN(\REGF/pbmemout1/n5913 ), .A(
        \pk_s89l_h[7] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[7] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[7] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[7] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U445  ( .ZN(\REGF/pbmemout1/n6066 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(1'b0), .F(
        \pk_rread_h[6] ), .G(\REGF/pk_idcz_h[27] ), .H(\pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U837  ( .ZN(\REGF/pbmemout1/n6380 ), .A(
        \pk_sra1_h[0] ), .B(\pk_rread_h[44] ), .C(CDOUT[0]), .D(
        \pk_rread_h[45] ), .E(CDOUT[32]), .F(\pk_rread_h[46] ), .G(1'b0), .H(
        \pk_rread_h[47] ) );
    snl_nand04x0 \REGF/pbmemout1/U268  ( .ZN(\REGF/pbmemout1/n5771 ), .A(
        \REGF/pbmemout1/n5924 ), .B(\REGF/pbmemout1/n5923 ), .C(
        \REGF/pbmemout1/n5922 ), .D(\REGF/pbmemout1/n5921 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U749  ( .ZN(\REGF/pbmemout1/n6309 ), .A(
        \pk_scba_h[13] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[13] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[13] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[13] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U479  ( .ZN(\REGF/pbmemout1/n6093 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \pk_stat_h[0] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] )
         );
    snl_oai022x1 \REGF/pbmemout1/U44  ( .ZN(\pk_ada_h[0] ), .A(
        \REGF/pbmemout1/n5677 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5679 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U56  ( .ZN(\pk_ada_h[12] ), .A(
        \REGF/pbmemout1/n5703 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5704 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_oai022x1 \REGF/pbmemout1/U94  ( .ZN(\REGF/pbmemout1/O_LDO[18] ), .A(
        \REGF/pbmemout1/n5715 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5716 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U136  ( .Z(\pk_pdo_h[28] ), .A(
        \REGF/pbmemout1/n5857 ), .B(\REGF/pbmemout1/n5858 ), .C(
        \REGF/pbmemout1/n5859 ), .D(\REGF/pbmemout1/n5860 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U354  ( .ZN(\REGF/pbmemout1/n5993 ), .A(
        \pk_s89l_h[31] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[31] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[31] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[31] ), .H(\pk_rread_h[35] ) );
    snl_nand04x0 \REGF/pbmemout1/U373  ( .ZN(\REGF/pbmemout1/n5868 ), .A(
        \REGF/pbmemout1/n6008 ), .B(\REGF/pbmemout1/n6007 ), .C(
        \REGF/pbmemout1/n6006 ), .D(\REGF/pbmemout1/n6005 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U545  ( .ZN(\REGF/pbmemout1/n6146 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[22] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[22] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U562  ( .ZN(\REGF/pbmemout1/n6160 ), .A(
        \pk_spr_h[22] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[22] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[22] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[22] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U652  ( .ZN(\REGF/pbmemout1/n6232 ), .A(
        \REGF/pk_s0ba_h[18] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[18] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[18] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[18] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U675  ( .ZN(\REGF/pbmemout1/n6250 ), .A(
        \pk_s01l_h[17] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[13] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[17] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[17] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U727  ( .ZN(\REGF/pbmemout1/n6292 ), .A(
        \pk_pcs1_h[14] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[14] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[14] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[14] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U206  ( .ZN(\REGF/pbmemout1/n5875 ), .A(
        \pk_rread_h[8] ), .B(\pk_idcy_h[9] ), .C(\pk_rread_h[9] ), .D(
        \pk_idcx_h[9] ), .E(\pk_rread_h[10] ), .F(\pk_idcw_h[9] ), .G(
        \pk_rread_h[11] ), .H(\pk_pcs2_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U396  ( .ZN(\REGF/pbmemout1/n6027 ), .A(1'b0
        ), .B(\pk_rread_h[40] ), .C(\pk_psae_h[2] ), .D(\pk_rread_h[41] ), .E(
        \REGF/RO_SRDA[2] ), .F(\pk_rread_h[42] ), .G(\pk_sra2_h[2] ), .H(
        \pk_rread_h[43] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U417  ( .ZN(\REGF/pbmemout1/n6044 ), .A(
        \pk_sra1_h[29] ), .B(\pk_rread_h[44] ), .C(CDOUT[29]), .D(
        \pk_rread_h[45] ), .E(1'b0), .F(\pk_rread_h[46] ), .G(CDOUT[57]), .H(
        \pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U587  ( .ZN(\REGF/pbmemout1/n6180 ), .A(1'b0
        ), .B(\pk_rread_h[12] ), .C(1'b0), .D(\pk_rread_h[13] ), .E(1'b0), .F(
        \pk_rread_h[14] ), .G(1'b0), .H(\pk_rread_h[15] ) );
    snl_oai022x1 \REGF/pbmemout1/U71  ( .ZN(\pk_ada_h[27] ), .A(
        \REGF/pbmemout1/n5733 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5734 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U221  ( .ZN(\REGF/pbmemout1/n5887 ), .A(
        \pk_rread_h[56] ), .B(\pk_indz_h[9] ), .C(\pk_rread_h[57] ), .D(
        \pk_indy_h[9] ), .E(\pk_rread_h[58] ), .F(\pk_indx_h[9] ), .G(
        \pk_rread_h[59] ), .H(\pk_indw_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U842  ( .ZN(\REGF/pbmemout1/n6384 ), .A(
        \pk_spr_h[0] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[0] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[0] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[0] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U430  ( .ZN(\REGF/pbmemout1/n6054 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_or04x1 \REGF/pbmemout1/U111  ( .Z(\pk_pdo_h[3] ), .A(
        \REGF/pbmemout1/n5757 ), .B(\REGF/pbmemout1/n5758 ), .C(
        \REGF/pbmemout1/n5759 ), .D(\REGF/pbmemout1/n5760 ) );
    snl_or04x1 \REGF/pbmemout1/U124  ( .Z(\pk_pdo_h[16] ), .A(
        \REGF/pbmemout1/n5809 ), .B(\REGF/pbmemout1/n5810 ), .C(
        \REGF/pbmemout1/n5811 ), .D(\REGF/pbmemout1/n5812 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U690  ( .ZN(\REGF/pbmemout1/n6262 ), .A(
        \pk_s8ba_h[16] ), .B(\pk_rread_h[20] ), .C(\pk_s7ba_h[16] ), .D(
        \pk_rread_h[21] ), .E(\pk_s6ba_h[16] ), .F(\pk_rread_h[22] ), .G(
        \pk_s5ba_h[16] ), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U700  ( .ZN(\REGF/pbmemout1/n6270 ), .A(
        \REGF/RO_PCON[16] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[16] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[16] ), .F(\pk_rread_h[54] ), .G(
        \REGF/pk_stat_h[16] ), .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U214  ( .ZN(\REGF/pbmemout1/n5881 ), .A(
        \pk_rread_h[32] ), .B(\pk_s89l_h[9] ), .C(\pk_rread_h[33] ), .D(
        \pk_s67l_h[9] ), .E(\pk_rread_h[34] ), .F(\pk_s45l_h[9] ), .G(
        \pk_rread_h[35] ), .H(\pk_s23l_h[9] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U595  ( .ZN(\REGF/pbmemout1/n6186 ), .A(
        \pk_s01l_h[20] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[16] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[20] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[20] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U735  ( .ZN(\REGF/pbmemout1/n6298 ), .A(
        \pk_s01l_h[14] ), .B(\pk_rread_h[36] ), .C(1'b0), .D(\pk_rread_h[37] ), 
        .E(\pk_trba_h[14] ), .F(\pk_rread_h[38] ), .G(\REGF/RO_ERRA[14] ), .H(
        \pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U384  ( .ZN(\REGF/pbmemout1/n6017 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(\REGF/pk_exco_h[2] ), .D(\pk_rread_h[1] ), 
        .E(\REGF/pk_scti_h[2] ), .F(\pk_rread_h[2] ), .G(\pk_sati_h[2] ), .H(
        \pk_rread_h[3] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U405  ( .ZN(\REGF/pbmemout1/n6034 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_hh[29] ), .F(\pk_rread_h[6] ), .G(\REGF/pk_idcz_h[29] ), .H(
        \pk_rread_h[7] ) );
    snl_oai022x1 \REGF/pbmemout1/U63  ( .ZN(\pk_ada_h[19] ), .A(
        \REGF/pbmemout1/n5717 ), .B(\REGF/pbmemout1/n5678 ), .C(
        \REGF/pbmemout1/n5718 ), .D(\REGF/pbmemout1/n5680 ) );
    snl_nand04x0 \REGF/pbmemout1/U233  ( .ZN(\REGF/pbmemout1/n5780 ), .A(
        \REGF/pbmemout1/n5896 ), .B(\REGF/pbmemout1/n5895 ), .C(
        \REGF/pbmemout1/n5894 ), .D(\REGF/pbmemout1/n5893 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U422  ( .ZN(\REGF/pbmemout1/n6048 ), .A(
        \pk_spr_h[29] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[29] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[29] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[29] ), .H(\pk_rread_h[63] ) );
    snl_oai022x1 \REGF/pbmemout1/U86  ( .ZN(\REGF/pbmemout1/O_LDO[10] ), .A(
        \REGF/pbmemout1/n5699 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5700 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_oai022x1 \REGF/pbmemout1/U103  ( .ZN(\REGF/pbmemout1/O_LDO[27] ), .A(
        \REGF/pbmemout1/n5733 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5734 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U712  ( .ZN(\REGF/pbmemout1/n6280 ), .A(
        \pk_s0ba_h[15] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[15] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[15] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[15] ), .H(\pk_rread_h[31] ) );
    snl_invx05 \REGF/pbmemout1/U188  ( .ZN(\REGF/pbmemout1/n5712 ), .A(
        \REGF/RO_EACC[16] ) );
    snl_nand04x0 \REGF/pbmemout1/U328  ( .ZN(\REGF/pbmemout1/n5759 ), .A(
        \REGF/pbmemout1/n5972 ), .B(\REGF/pbmemout1/n5971 ), .C(
        \REGF/pbmemout1/n5970 ), .D(\REGF/pbmemout1/n5969 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U682  ( .ZN(\REGF/pbmemout1/n6256 ), .A(
        \pk_spr_h[17] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[17] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[17] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[17] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U539  ( .ZN(\REGF/pbmemout1/n6141 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \pk_stat_h[18] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] )
         );
    snl_aoi2222x0 \REGF/pbmemout1/U799  ( .ZN(\REGF/pbmemout1/n6349 ), .A(
        ph_izco_h), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        CDOUT[41]), .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U609  ( .ZN(\REGF/pbmemout1/n6197 ), .A(
        \pk_scba_h[1] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[1] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[1] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[1] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U346  ( .ZN(\REGF/pbmemout1/n5987 ), .A(
        \REGF/pk_idcy_h[31] ), .B(\pk_rread_h[8] ), .C(\REGF/pk_idcx_h[31] ), 
        .D(\pk_rread_h[9] ), .E(\REGF/pk_idcw_h[31] ), .F(\pk_rread_h[10] ), 
        .G(1'b0), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U557  ( .ZN(\REGF/pbmemout1/n6156 ), .A(
        \pk_sra1_h[22] ), .B(\pk_rread_h[44] ), .C(CDOUT[22]), .D(
        \pk_rread_h[45] ), .E(CDOUT[54]), .F(\pk_rread_h[46] ), .G(
        \REGF/RO_PSTA[22] ), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U361  ( .ZN(\REGF/pbmemout1/n5999 ), .A(
        \REGF/pk_indz_h[31] ), .B(\pk_rread_h[56] ), .C(\REGF/pk_indy_h[31] ), 
        .D(\pk_rread_h[57] ), .E(\REGF/pk_indx_h[31] ), .F(\pk_rread_h[58] ), 
        .G(\REGF/pk_indw_h[31] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U640  ( .ZN(\REGF/pbmemout1/n6222 ), .A(
        \REGF/RO_PCON[19] ), .B(\pk_rread_h[52] ), .C(1'b0), .D(
        \pk_rread_h[53] ), .E(1'b0), .F(\pk_rread_h[54] ), .G(1'b0), .H(
        \pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U667  ( .ZN(\REGF/pbmemout1/n6244 ), .A(
        \pk_pcs1_h[17] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[17] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[17] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[17] ), .H(\pk_rread_h[15] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U570  ( .ZN(\REGF/pbmemout1/n6166 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U819  ( .ZN(\REGF/pbmemout1/n6365 ), .A(
        ph_iyco_h), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        CDOUT[40]), .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_invx05 \REGF/pbmemout1/U151  ( .ZN(\REGF/pbmemout1/n5687 ), .A(
        \REGF/RO_ACC[4] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U261  ( .ZN(\REGF/pbmemout1/n5919 ), .A(
        \pk_indz_h[7] ), .B(\pk_rread_h[56] ), .C(\pk_indy_h[7] ), .D(
        \pk_rread_h[57] ), .E(\pk_indx_h[7] ), .F(\pk_rread_h[58] ), .G(
        \pk_indw_h[7] ), .H(\pk_rread_h[59] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U470  ( .ZN(\REGF/pbmemout1/n6086 ), .A(1'b0
        ), .B(\pk_rread_h[20] ), .C(1'b0), .D(\pk_rread_h[21] ), .E(1'b0), .F(
        \pk_rread_h[22] ), .G(1'b0), .H(\pk_rread_h[23] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U740  ( .ZN(\REGF/pbmemout1/n6302 ), .A(
        \REGF/RO_PCON[14] ), .B(\pk_rread_h[52] ), .C(\REGF/RO_PPCN[14] ), .D(
        \pk_rread_h[53] ), .E(\pk_pc_h[14] ), .F(\pk_rread_h[54] ), .G(1'b0), 
        .H(\pk_rread_h[55] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U802  ( .ZN(\REGF/pbmemout1/n6352 ), .A(
        \pk_spr_h[11] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[11] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[11] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[11] ), .H(\pk_rread_h[63] ) );
    snl_invx05 \REGF/pbmemout1/U176  ( .ZN(\REGF/pbmemout1/n5722 ), .A(
        \REGF/RO_EACC[21] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U767  ( .ZN(\REGF/pbmemout1/n6324 ), .A(
        \pk_pcs1_h[12] ), .B(\pk_rread_h[12] ), .C(\pk_sfba_h[12] ), .D(
        \pk_rread_h[13] ), .E(\pk_seba_h[12] ), .F(\pk_rread_h[14] ), .G(
        \pk_sdba_h[12] ), .H(\pk_rread_h[15] ) );
    snl_oai022x1 \REGF/pbmemout1/U78  ( .ZN(\REGF/pbmemout1/O_LDO[2] ), .A(
        \REGF/pbmemout1/n5683 ), .B(\REGF/pbmemout1/n5743 ), .C(
        \REGF/pbmemout1/n5684 ), .D(\REGF/pbmemout1/n5744 ) );
    snl_or04x1 \REGF/pbmemout1/U118  ( .Z(\pk_pdo_h[10] ), .A(
        \REGF/pbmemout1/n5785 ), .B(\REGF/pbmemout1/n5786 ), .C(
        \REGF/pbmemout1/n5787 ), .D(\REGF/pbmemout1/n5788 ) );
    snl_invx05 \REGF/pbmemout1/U193  ( .ZN(\REGF/pbmemout1/n5707 ), .A(
        \REGF/RO_ACC[14] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U246  ( .ZN(\REGF/pbmemout1/n5907 ), .A(
        \pk_idcy_h[7] ), .B(\pk_rread_h[8] ), .C(\pk_idcx_h[7] ), .D(
        \pk_rread_h[9] ), .E(\pk_idcw_h[7] ), .F(\pk_rread_h[10] ), .G(
        \pk_pcs2_h[7] ), .H(\pk_rread_h[11] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U457  ( .ZN(\REGF/pbmemout1/n6076 ), .A(1'b0
        ), .B(\pk_rread_h[44] ), .C(CDOUT[27]), .D(\pk_rread_h[45] ), .E(CDOUT
        [59]), .F(\pk_rread_h[46] ), .G(CDOUT[55]), .H(\pk_rread_h[47] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U782  ( .ZN(\REGF/pbmemout1/n6336 ), .A(
        \pk_spr_h[12] ), .B(\pk_rread_h[60] ), .C(\pk_dpr_h[12] ), .D(
        \pk_rread_h[61] ), .E(\REGF/RO_EACC[12] ), .F(\pk_rread_h[62] ), .G(
        \REGF/RO_ACC[12] ), .H(\pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U825  ( .ZN(\REGF/pbmemout1/n6370 ), .A(
        pk_sased_h), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(
        \pk_saco_lh[0] ), .F(\pk_rread_h[6] ), .G(\pk_idcz_h[0] ), .H(
        \pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U284  ( .ZN(\REGF/pbmemout1/n5937 ), .A(1'b0
        ), .B(\pk_rread_h[0] ), .C(1'b0), .D(\pk_rread_h[1] ), .E(
        \REGF/pk_scti_h[5] ), .F(\pk_rread_h[2] ), .G(1'b0), .H(
        \pk_rread_h[3] ) );
    snl_nand04x0 \REGF/pbmemout1/U333  ( .ZN(\REGF/pbmemout1/n5760 ), .A(
        \REGF/pbmemout1/n5976 ), .B(\REGF/pbmemout1/n5975 ), .C(
        \REGF/pbmemout1/n5974 ), .D(\REGF/pbmemout1/n5973 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U612  ( .ZN(\REGF/pbmemout1/n6200 ), .A(
        \pk_s0ba_h[1] ), .B(\pk_rread_h[28] ), .C(\pk_sefl_h[1] ), .D(
        \pk_rread_h[29] ), .E(\pk_scdl_h[1] ), .F(\pk_rread_h[30] ), .G(
        \pk_sabl_h[1] ), .H(\pk_rread_h[31] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U505  ( .ZN(\REGF/pbmemout1/n6114 ), .A(1'b0
        ), .B(\pk_rread_h[4] ), .C(1'b0), .D(\pk_rread_h[5] ), .E(1'b0), .F(
        \pk_rread_h[6] ), .G(\REGF/pk_idcz_h[24] ), .H(\pk_rread_h[7] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U522  ( .ZN(\REGF/pbmemout1/n6128 ), .A(1'b0
        ), .B(\pk_rread_h[60] ), .C(1'b0), .D(\pk_rread_h[61] ), .E(
        \REGF/RO_EACC[24] ), .F(\pk_rread_h[62] ), .G(\REGF/RO_ACC[24] ), .H(
        \pk_rread_h[63] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U314  ( .ZN(\REGF/pbmemout1/n5961 ), .A(
        \pk_s89l_h[4] ), .B(\pk_rread_h[32] ), .C(\pk_s67l_h[4] ), .D(
        \pk_rread_h[33] ), .E(\pk_s45l_h[4] ), .F(\pk_rread_h[34] ), .G(
        \pk_s23l_h[4] ), .H(\pk_rread_h[35] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U495  ( .ZN(\REGF/pbmemout1/n6106 ), .A(
        \pk_s01l_h[25] ), .B(\pk_rread_h[36] ), .C(\REGF/RO_TRCO[25] ), .D(
        \pk_rread_h[37] ), .E(1'b0), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[25] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U635  ( .ZN(\REGF/pbmemout1/n6218 ), .A(
        \pk_s01l_h[19] ), .B(\pk_rread_h[36] ), .C(\pk_stdat[15] ), .D(
        \pk_rread_h[37] ), .E(\pk_trba_h[19] ), .F(\pk_rread_h[38] ), .G(
        \REGF/RO_ERRA[19] ), .H(\pk_rread_h[39] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U709  ( .ZN(\REGF/pbmemout1/n6277 ), .A(
        \pk_scba_h[15] ), .B(\pk_rread_h[16] ), .C(\pk_sbba_h[15] ), .D(
        \pk_rread_h[17] ), .E(\pk_saba_h[15] ), .F(\pk_rread_h[18] ), .G(
        \pk_s9ba_h[15] ), .H(\pk_rread_h[19] ) );
    snl_aoi2222x0 \REGF/pbmemout1/U699  ( .ZN(\REGF/pbmemout1/n6269 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(
        \REGF/RO_PSTA[16] ), .F(\pk_rread_h[50] ), .G(1'b0), .H(
        \pk_rread_h[51] ) );
    snl_nand04x0 \REGF/pbmemout1/U228  ( .ZN(\REGF/pbmemout1/n5779 ), .A(
        \REGF/pbmemout1/n5892 ), .B(\REGF/pbmemout1/n5891 ), .C(
        \REGF/pbmemout1/n5890 ), .D(\REGF/pbmemout1/n5889 ) );
    snl_aoi2222x0 \REGF/pbmemout1/U439  ( .ZN(\REGF/pbmemout1/n6061 ), .A(1'b0
        ), .B(\pk_rread_h[48] ), .C(1'b0), .D(\pk_rread_h[49] ), .E(CDOUT[56]), 
        .F(\pk_rread_h[50] ), .G(1'b0), .H(\pk_rread_h[51] ) );
    snl_nand12x8 \REGF/pbmemff11/U619  ( .ZN(\REGF/pbmemff11/n_1556 ), .A(
        \pk_rwrit_h[66] ), .B(\REGF/pbmemff11/n5643 ) );
    snl_and02x1 \REGF/pbmemff11/U692  ( .Z(\REGF/pbmemff11/RO_ACC147[29] ), 
        .A(\REGF/RI_ACC[29] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U840  ( .ZN(\REGF/pbmemff11/RO_INDX349[21] ), 
        .A(\REGF/pbmemff11/n5125 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[8]  ( .Q(\REGF/RO_EACC[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_EACC187[8] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U702  ( .ZN(\REGF/pbmemff11/RO_INDW309[7] ), 
        .A(\REGF/pbmemff11/n5111 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U725  ( .ZN(\REGF/pbmemff11/RO_INDW309[30] ), 
        .A(\REGF/pbmemff11/n5134 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[25]  ( .Q(\REGF/pk_indx_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[25] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U867  ( .ZN(\REGF/pbmemff11/RO_INDZ429[16] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5120 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[16]  ( .Q(\pk_indx_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[16] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[3]  ( .Q(\pk_dpr_h[3] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[3] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U625  ( .Z(\REGF/pbmemff11/n5096 ), .A(
        \REGF/pbmemff11/n5100 ), .B(\REGF/pbmemff11/n5643 ) );
    snl_nand12x1 \REGF/pbmemff11/U650  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[15] 
        ), .A(\REGF/RI_DPR[15] ), .B(\pk_rwrit_h[66] ) );
    snl_nor02x1 \REGF/pbmemff11/U789  ( .ZN(\REGF/pbmemff11/RO_INDY389[2] ), 
        .A(\REGF/pbmemff11/n5106 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[1]  ( .Q(\pk_indx_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDX349[1] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_and02x1 \REGF/pbmemff11/U677  ( .Z(\REGF/pbmemff11/RO_ACC147[14] ), 
        .A(\REGF/RI_ACC[14] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U882  ( .ZN(\REGF/pbmemff11/RO_INDZ429[31] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5135 ) );
    snl_invx05 \REGF/pbmemff11/U912  ( .ZN(\REGF/pbmemff11/n5122 ), .A(PDLIN
        [18]) );
    snl_and02x1 \REGF/pbmemff11/U750  ( .Z(\REGF/pbmemff11/RO_EACC187[23] ), 
        .A(\REGF/RI_EACC[23] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U777  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[18] 
        ), .A(\REGF/RI_SPR[18] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U809  ( .ZN(\REGF/pbmemff11/RO_INDY389[22] ), 
        .A(\REGF/pbmemff11/n5126 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[6]  ( .Q(\pk_indy_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDY389[6] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[3]  ( .Q(\pk_indw_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[3] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_STAT5B_reg[5]  ( .Q(\REGF/pk_stat_h[31] 
        ), .D(1'b0), .EN(\REGF/pbmemff11/n5643 ), .RN(\REGF/pbmemff11/n5091 ), 
        .SD(\REGF/RI_STAT[5] ), .SE(\pk_rwrit_h[60] ), .CP(SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U812  ( .ZN(\REGF/pbmemff11/RO_INDY389[25] ), 
        .A(\REGF/pbmemff11/n5129 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U835  ( .ZN(\REGF/pbmemff11/RO_INDX349[16] ), 
        .A(\REGF/pbmemff11/n5120 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_invx05 \REGF/pbmemff11/U899  ( .ZN(\REGF/pbmemff11/n5106 ), .A(PDLIN
        [2]) );
    snl_invx05 \REGF/pbmemff11/U909  ( .ZN(\REGF/pbmemff11/n5124 ), .A(PDLIN
        [20]) );
    snl_and02x1 \REGF/pbmemff11/U689  ( .Z(\REGF/pbmemff11/RO_ACC147[26] ), 
        .A(\REGF/RI_ACC[26] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U792  ( .ZN(\REGF/pbmemff11/RO_INDY389[5] ), 
        .A(\REGF/pbmemff11/n5109 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[1]  ( .Q(\REGF/RO_EACC[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[1] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[3]  ( .Q(\REGF/RO_ACC[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_ACC147[3] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_nor02x1 \REGF/pbmemff11/U719  ( .ZN(\REGF/pbmemff11/RO_INDW309[24] ), 
        .A(\REGF/pbmemff11/n5128 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[7]  ( .Q(\pk_indw_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[7] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[8]  ( .Q(\pk_indx_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDX349[8] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_ffqrnx1 \REGF/pbmemff11/RO_STAT5B_reg[1]  ( .Q(\pk_stat_h[1] ), .D(
        \REGF/pbmemff11/RO_STAT5BP[1] ), .RN(\REGF/pbmemff11/n5091 ), .CP(SCLK
        ) );
    snl_invx2 \REGF/pbmemff11/U611  ( .ZN(\REGF/pbmemff11/n5093 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_invx2 \REGF/pbmemff11/U616  ( .ZN(\REGF/pbmemff11/n5091 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_invx2 \REGF/pbmemff11/U617  ( .ZN(\REGF/pbmemff11/n5090 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_nand12x1 \REGF/pbmemff11/U637  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[2] ), 
        .A(\REGF/RI_DPR[2] ), .B(\pk_rwrit_h[66] ) );
    snl_nor02x1 \REGF/pbmemff11/U849  ( .ZN(\REGF/pbmemff11/RO_INDX349[30] ), 
        .A(\REGF/pbmemff11/n5134 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[2]  ( .Q(\pk_indy_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDY389[2] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_nand12x1 \REGF/pbmemff11/U642  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[7] ), 
        .A(\REGF/RI_DPR[7] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U659  ( .Z(\REGF/pbmemff11/RO_DPR28B227[24] ), 
        .A(\REGF/RI_DPR[24] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U780  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[21] 
        ), .A(\REGF/RI_SPR[21] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[5]  ( .Q(\pk_indx_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDX349[5] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_and02x1 \REGF/pbmemff11/U742  ( .Z(\REGF/pbmemff11/RO_EACC187[15] ), 
        .A(\REGF/RI_EACC[15] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U765  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[6] ), 
        .A(\REGF/RI_SPR[6] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U800  ( .ZN(\REGF/pbmemff11/RO_INDY389[13] ), 
        .A(\REGF/pbmemff11/n5117 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U827  ( .ZN(\REGF/pbmemff11/RO_INDX349[8] ), 
        .A(\REGF/pbmemff11/n5112 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[21]  ( .Q(\pk_indx_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[21] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[12]  ( .Q(\pk_indx_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDX349[12] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[7]  ( .Q(\pk_dpr_h[7] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[7] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U759  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[0] ), 
        .A(\REGF/RI_SPR[0] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[7]  ( .Q(\REGF/RO_ACC[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_ACC147[7] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_nand12x1 \REGF/pbmemff11/U645  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[10] 
        ), .A(\REGF/RI_DPR[10] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U662  ( .Z(\REGF/pbmemff11/RO_DPR28B227[27] ), 
        .A(\REGF/RI_DPR[27] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U665  ( .Z(\REGF/pbmemff11/RO_ACC147[2] ), .A(
        \REGF/RI_ACC[2] ), .B(\pk_rwrit_h[68] ) );
    snl_invx05 \REGF/pbmemff11/U890  ( .ZN(\REGF/pbmemff11/n5113 ), .A(PDLIN
        [9]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[5]  ( .Q(\REGF/RO_EACC[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_EACC187[5] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U900  ( .ZN(\REGF/pbmemff11/n5133 ), .A(PDLIN
        [29]) );
    snl_nand02x1 \REGF/pbmemff11/U927  ( .ZN(\REGF/pbmemff11/n5138 ), .A(
        \REGF/pbmemff11/n5145 ), .B(\REGF/pbmemff11/n5137 ) );
    snl_and02x1 \REGF/pbmemff11/U680  ( .Z(\REGF/pbmemff11/RO_ACC147[17] ), 
        .A(\REGF/RI_ACC[17] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U710  ( .ZN(\REGF/pbmemff11/RO_INDW309[15] ), 
        .A(\REGF/pbmemff11/n5119 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U852  ( .ZN(\REGF/pbmemff11/RO_INDZ429[1] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5105 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[31]  ( .Q(\REGF/pk_indx_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[31] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[28]  ( .Q(\REGF/pk_indx_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDX349[28] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U687  ( .Z(\REGF/pbmemff11/RO_ACC147[24] ), 
        .A(\REGF/RI_ACC[24] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U730  ( .Z(\REGF/pbmemff11/RO_EACC187[3] ), 
        .A(\REGF/RI_EACC[3] ), .B(\pk_rwrit_h[67] ) );
    snl_and02x1 \REGF/pbmemff11/U737  ( .Z(\REGF/pbmemff11/RO_EACC187[10] ), 
        .A(\REGF/RI_EACC[10] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U872  ( .ZN(\REGF/pbmemff11/RO_INDZ429[21] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5125 ) );
    snl_nor02x1 \REGF/pbmemff11/U875  ( .ZN(\REGF/pbmemff11/RO_INDZ429[24] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5128 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[9]  ( .Q(\pk_indy_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDY389[9] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_nor02x1 \REGF/pbmemff11/U717  ( .ZN(\REGF/pbmemff11/RO_INDW309[22] ), 
        .A(\REGF/pbmemff11/n5126 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nand12x1 \REGF/pbmemff11/U779  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[20] 
        ), .A(\REGF/RI_SPR[20] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U855  ( .ZN(\REGF/pbmemff11/RO_INDZ429[4] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5108 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[5]  ( .Q(\REGF/RO_ACC[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_ACC147[5] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[7]  ( .Q(\REGF/RO_EACC[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[7] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U897  ( .ZN(\REGF/pbmemff11/n5135 ), .A(PDLIN
        [31]) );
    snl_invx05 \REGF/pbmemff11/U907  ( .ZN(\REGF/pbmemff11/n5126 ), .A(PDLIN
        [22]) );
    snl_invx05 \REGF/pbmemff11/U920  ( .ZN(\REGF/pbmemff11/n5114 ), .A(PDLIN
        [10]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[19]  ( .Q(\pk_indx_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDX349[19] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U679  ( .Z(\REGF/pbmemff11/RO_ACC147[16] ), 
        .A(\REGF/RI_ACC[16] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U745  ( .Z(\REGF/pbmemff11/RO_EACC187[18] ), 
        .A(\REGF/RI_EACC[18] ), .B(\pk_rwrit_h[67] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[23]  ( .Q(\pk_indx_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDX349[23] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[7]  ( .Q(\pk_indx_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[7] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_nand12x1 \REGF/pbmemff11/U762  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[3] ), 
        .A(\REGF/RI_SPR[3] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U807  ( .ZN(\REGF/pbmemff11/RO_INDY389[20] ), 
        .A(\REGF/pbmemff11/n5124 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[10]  ( .Q(\pk_indx_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[10] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[5]  ( .Q(\pk_dpr_h[5] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[5] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U820  ( .ZN(\REGF/pbmemff11/RO_INDX349[1] ), 
        .A(\REGF/pbmemff11/n5105 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U869  ( .ZN(\REGF/pbmemff11/RO_INDZ429[18] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5122 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[5]  ( .Q(\pk_indw_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[5] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[0]  ( .Q(\pk_indy_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[0] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_ffqrnx1 \REGF/pbmemff11/RO_STAT5B_reg[3]  ( .Q(\pk_stat_h[18] ), .D(
        \REGF/pbmemff11/RO_STAT5BP[3] ), .RN(\REGF/pbmemff11/n5091 ), .CP(SCLK
        ) );
    snl_nand12x8 \REGF/pbmemff11/U622  ( .ZN(\REGF/pbmemff11/n_1032 ), .A(
        \pk_rwrit_h[67] ), .B(\REGF/pbmemff11/n5643 ) );
    snl_invx1 \REGF/pbmemff11/U630  ( .ZN(\REGF/pbmemff11/n5100 ), .A(
        \pk_rwrit_h[64] ) );
    snl_nor02x1 \REGF/pbmemff11/U787  ( .ZN(\REGF/pbmemff11/RO_INDY389[0] ), 
        .A(\REGF/pbmemff11/n5104 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U795  ( .ZN(\REGF/pbmemff11/RO_INDY389[8] ), 
        .A(\REGF/pbmemff11/n5112 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[8]  ( .Q(\pk_dpr_h[8] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[8] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U639  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[4] ), 
        .A(\REGF/RI_DPR[4] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U657  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[22] 
        ), .A(\REGF/RI_DPR[22] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U670  ( .Z(\REGF/pbmemff11/RO_ACC147[7] ), .A(
        \REGF/RI_ACC[7] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U739  ( .Z(\REGF/pbmemff11/RO_EACC187[12] ), 
        .A(\REGF/RI_EACC[12] ), .B(\pk_rwrit_h[67] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[1]  ( .Q(\REGF/RO_ACC[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_ACC147[1] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[3]  ( .Q(\REGF/RO_EACC[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[3] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U757  ( .Z(\REGF/pbmemff11/RO_EACC187[30] ), 
        .A(\REGF/RI_EACC[30] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U770  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[11] 
        ), .A(\REGF/RI_SPR[11] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U815  ( .ZN(\REGF/pbmemff11/RO_INDY389[28] ), 
        .A(\REGF/pbmemff11/n5132 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U832  ( .ZN(\REGF/pbmemff11/RO_INDX349[13] ), 
        .A(\REGF/pbmemff11/n5117 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_muxi21x1 \REGF/pbmemff11/U929  ( .ZN(\REGF/pbmemff11/n5139 ), .A(
        \REGF/RI_STAT[2] ), .B(\REGF/pk_stat_h[16] ), .S(
        \REGF/pbmemff11/n5144 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[8]  ( .Q(\pk_indw_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[8] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_ao023x1 \REGF/pbmemff11/U885  ( .Z(\REGF/pbmemff11/RO_STAT5BP[1] ), 
        .A(\REGF/pbmemff11/n5136 ), .B(\REGF/pbmemff11/n5140 ), .C(
        \pk_stat_h[1] ), .D(\REGF/RI_STAT[1] ), .E(\REGF/pbmemff11/n5141 ) );
    snl_invx05 \REGF/pbmemff11/U915  ( .ZN(\REGF/pbmemff11/n5119 ), .A(PDLIN
        [15]) );
    snl_nor02x1 \REGF/pbmemff11/U695  ( .ZN(\REGF/pbmemff11/RO_INDW309[0] ), 
        .A(\REGF/pbmemff11/n5104 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U705  ( .ZN(\REGF/pbmemff11/RO_INDW309[10] ), 
        .A(\REGF/pbmemff11/n5114 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U722  ( .ZN(\REGF/pbmemff11/RO_INDW309[27] ), 
        .A(\REGF/pbmemff11/n5131 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U829  ( .ZN(\REGF/pbmemff11/RO_INDX349[10] ), 
        .A(\REGF/pbmemff11/n5114 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[4]  ( .Q(\pk_indy_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[4] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_nor02x1 \REGF/pbmemff11/U860  ( .ZN(\REGF/pbmemff11/RO_INDZ429[9] ), 
        .A(\REGF/pbmemff11/n5113 ), .B(\REGF/pbmemff11/n5103 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[1]  ( .Q(\pk_indw_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[1] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_nor02x1 \REGF/pbmemff11/U847  ( .ZN(\REGF/pbmemff11/RO_INDX349[28] ), 
        .A(\REGF/pbmemff11/n5132 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[27]  ( .Q(\REGF/pk_indx_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[27] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[14]  ( .Q(\pk_indx_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDX349[14] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[1]  ( .Q(\pk_dpr_h[1] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[1] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[3]  ( .Q(\pk_indx_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[3] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_and02x1 \REGF/pbmemff11/U786  ( .Z(\REGF/pbmemff11/RO_SPR28B268[27] ), 
        .A(\REGF/RI_SPR[27] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U868  ( .ZN(\REGF/pbmemff11/RO_INDZ429[17] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5121 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[8]  ( .Q(\REGF/RO_ACC[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_ACC147[8] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_invx1 \REGF/pbmemff11/U618  ( .ZN(\REGF/pbmemff11/n5089 ), .A(
        \REGF/n8052 ) );
    snl_bufx1 \REGF/pbmemff11/U623  ( .Z(\REGF/pbmemff11/n5094 ), .A(
        \REGF/pbmemff11/n_4044 ) );
    snl_invx1 \REGF/pbmemff11/U631  ( .ZN(\REGF/pbmemff11/n5102 ), .A(
        \pk_rwrit_h[62] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[17]  ( .Q(\pk_indy_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[17] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U638  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[3] ), 
        .A(\REGF/RI_DPR[3] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U644  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[9] ), 
        .A(\REGF/RI_DPR[9] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U663  ( .Z(\REGF/pbmemff11/RO_ACC147[0] ), .A(
        \REGF/RI_ACC[0] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U678  ( .Z(\REGF/pbmemff11/RO_ACC147[15] ), 
        .A(\REGF/RI_ACC[15] ), .B(\pk_rwrit_h[68] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[30]  ( .Q(\REGF/RO_ACC[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_ACC147[30] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[29]  ( .Q(\REGF/RO_ACC[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_ACC147[29] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[24]  ( .Q(\REGF/pk_indy_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDY389[24] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[16]  ( .Q(\pk_indz_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[16] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[18]  ( .Q(\pk_spr_h[18] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[18] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U744  ( .Z(\REGF/pbmemff11/RO_EACC187[17] ), 
        .A(\REGF/RI_EACC[17] ), .B(\pk_rwrit_h[67] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[25]  ( .Q(\REGF/pk_indz_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[25] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U763  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[4] ), 
        .A(\REGF/RI_SPR[4] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U806  ( .ZN(\REGF/pbmemff11/RO_INDY389[19] ), 
        .A(\REGF/pbmemff11/n5123 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[27]  ( .Q(\REGF/RO_EACC[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[27] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U821  ( .ZN(\REGF/pbmemff11/RO_INDX349[2] ), 
        .A(\REGF/pbmemff11/n5106 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[14]  ( .Q(\REGF/RO_EACC[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[14] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U778  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[19] 
        ), .A(\REGF/RI_SPR[19] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[20]  ( .Q(\REGF/RO_ACC[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_ACC147[20] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[13]  ( .Q(\REGF/RO_ACC[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_ACC147[13] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[7]  ( .Q(\pk_indz_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[7] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[22]  ( .Q(\pk_spr_h[22] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[22] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[11]  ( .Q(\pk_spr_h[11] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[11] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U896  ( .ZN(\REGF/pbmemff11/n5107 ), .A(PDLIN
        [3]) );
    snl_invx05 \REGF/pbmemff11/U921  ( .ZN(\REGF/pbmemff11/n5104 ), .A(PDLIN
        [0]) );
    snl_invx05 \REGF/pbmemff11/U906  ( .ZN(\REGF/pbmemff11/n5127 ), .A(PDLIN
        [23]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[27]  ( .Q(\REGF/pk_indw_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[27] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U686  ( .Z(\REGF/pbmemff11/RO_ACC147[23] ), 
        .A(\REGF/RI_ACC[23] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U716  ( .ZN(\REGF/pbmemff11/RO_INDW309[21] ), 
        .A(\REGF/pbmemff11/n5125 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_and02x1 \REGF/pbmemff11/U731  ( .Z(\REGF/pbmemff11/RO_EACC187[4] ), 
        .A(\REGF/RI_EACC[4] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U873  ( .ZN(\REGF/pbmemff11/RO_INDZ429[22] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5126 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[14]  ( .Q(\pk_indw_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDW309[14] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[14]  ( .Q(\pk_dpr_h[14] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[14] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_DPR28B_reg[27]  ( .Q(\pk_dpr_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[27] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U694  ( .Z(\REGF/pbmemff11/RO_ACC147[31] ), 
        .A(\REGF/RI_ACC[31] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U723  ( .ZN(\REGF/pbmemff11/RO_INDW309[28] ), 
        .A(\REGF/pbmemff11/n5132 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U854  ( .ZN(\REGF/pbmemff11/RO_INDZ429[3] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5107 ) );
    snl_nor02x1 \REGF/pbmemff11/U861  ( .ZN(\REGF/pbmemff11/RO_INDZ429[10] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5114 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[4]  ( .Q(\pk_spr_h[4] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[4] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[23]  ( .Q(\REGF/RO_EACC[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_EACC187[23] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[19]  ( .Q(\pk_indw_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[19] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U704  ( .ZN(\REGF/pbmemff11/RO_INDW309[9] ), 
        .A(\REGF/pbmemff11/n5113 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U846  ( .ZN(\REGF/pbmemff11/RO_INDX349[27] ), 
        .A(\REGF/pbmemff11/n5131 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[10]  ( .Q(\REGF/RO_EACC[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[10] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[21]  ( .Q(\pk_indz_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[21] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[12]  ( .Q(\pk_indz_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[12] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U656  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[21] 
        ), .A(\REGF/RI_DPR[21] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U671  ( .Z(\REGF/pbmemff11/RO_ACC147[8] ), .A(
        \REGF/RI_ACC[8] ), .B(\pk_rwrit_h[68] ) );
    snl_nand02x1 \REGF/pbmemff11/U884  ( .ZN(pk_ciffh), .A(
        \REGF/pbmemff11/n5139 ), .B(\REGF/pbmemff11/n5643 ) );
    snl_invx05 \REGF/pbmemff11/U914  ( .ZN(\REGF/pbmemff11/n5120 ), .A(PDLIN
        [16]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[20]  ( .Q(\pk_indy_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDY389[20] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[13]  ( .Q(\pk_indy_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDY389[13] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[9]  ( .Q(\pk_spr_h[9] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[9] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U756  ( .Z(\REGF/pbmemff11/RO_EACC187[29] ), 
        .A(\REGF/RI_EACC[29] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U828  ( .ZN(\REGF/pbmemff11/RO_INDX349[9] ), 
        .A(\REGF/pbmemff11/n5113 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[19]  ( .Q(\pk_dpr_h[19] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[19] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U771  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[12] 
        ), .A(\REGF/RI_SPR[12] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U814  ( .ZN(\REGF/pbmemff11/RO_INDY389[27] ), 
        .A(\REGF/pbmemff11/n5131 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[0]  ( .Q(\pk_spr_h[0] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[0] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U833  ( .ZN(\REGF/pbmemff11/RO_INDX349[14] ), 
        .A(\REGF/pbmemff11/n5118 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[30]  ( .Q(\REGF/pk_indy_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDY389[30] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[29]  ( .Q(\REGF/pk_indy_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[29] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U794  ( .ZN(\REGF/pbmemff11/RO_INDY389[7] ), 
        .A(\REGF/pbmemff11/n5111 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nand02x1 \REGF/pbmemff11/U928  ( .ZN(\REGF/pbmemff11/n5141 ), .A(
        \REGF/pbmemff11/n5145 ), .B(\REGF/pbmemff11/n5140 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[10]  ( .Q(\pk_dpr_h[10] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[10] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[19]  ( .Q(\REGF/RO_EACC[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[19] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[23]  ( .Q(\pk_dpr_h[23] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[23] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[23]  ( .Q(\pk_indw_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDW309[23] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[10]  ( .Q(\pk_indw_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[10] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_bufx1 \REGF/pbmemff11/U624  ( .Z(\REGF/pbmemff11/n5095 ), .A(
        \REGF/pbmemff11/n_3464 ) );
    snl_and02x1 \REGF/pbmemff11/U738  ( .Z(\REGF/pbmemff11/RO_EACC187[11] ), 
        .A(\REGF/RI_EACC[11] ), .B(\pk_rwrit_h[67] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[24]  ( .Q(\REGF/RO_ACC[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[24] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[17]  ( .Q(\REGF/RO_ACC[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[17] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_SPR28B_reg[26]  ( .Q(\pk_spr_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[26] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[3]  ( .Q(\pk_indz_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[3] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[15]  ( .Q(\pk_spr_h[15] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[15] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[31]  ( .Q(\REGF/pk_indz_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[31] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[28]  ( .Q(\REGF/pk_indz_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[28] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[21]  ( .Q(\pk_indw_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[21] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U651  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[16] 
        ), .A(\REGF/RI_DPR[16] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U688  ( .Z(\REGF/pbmemff11/RO_ACC147[25] ), 
        .A(\REGF/RI_ACC[25] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U718  ( .ZN(\REGF/pbmemff11/RO_INDW309[23] ), 
        .A(\REGF/pbmemff11/n5127 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U793  ( .ZN(\REGF/pbmemff11/RO_INDY389[6] ), 
        .A(\REGF/pbmemff11/n5110 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[31]  ( .Q(\REGF/RO_EACC[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_EACC187[31] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[28]  ( .Q(\REGF/RO_EACC[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_EACC187[28] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[12]  ( .Q(\pk_indw_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDW309[12] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[26]  ( .Q(\REGF/RO_ACC[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_ACC147[26] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[15]  ( .Q(\REGF/RO_ACC[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[15] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[1]  ( .Q(\pk_indz_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[1] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_SPR28B_reg[24]  ( .Q(\pk_spr_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[24] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[17]  ( .Q(\pk_spr_h[17] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[17] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U751  ( .Z(\REGF/pbmemff11/RO_EACC187[24] ), 
        .A(\REGF/RI_EACC[24] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U776  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[17] 
        ), .A(\REGF/RI_SPR[17] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[19]  ( .Q(\pk_indz_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[19] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U813  ( .ZN(\REGF/pbmemff11/RO_INDY389[26] ), 
        .A(\REGF/pbmemff11/n5130 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U834  ( .ZN(\REGF/pbmemff11/RO_INDX349[15] ), 
        .A(\REGF/pbmemff11/n5119 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[2]  ( .Q(\pk_spr_h[2] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[2] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[18]  ( .Q(\pk_indy_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDY389[18] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U898  ( .ZN(\REGF/pbmemff11/n5134 ), .A(PDLIN
        [30]) );
    snl_invx05 \REGF/pbmemff11/U908  ( .ZN(\REGF/pbmemff11/n5125 ), .A(PDLIN
        [21]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[11]  ( .Q(\pk_indy_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDY389[11] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[21]  ( .Q(\pk_dpr_h[21] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[21] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[12]  ( .Q(\pk_dpr_h[12] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[12] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U676  ( .Z(\REGF/pbmemff11/RO_ACC147[13] ), 
        .A(\REGF/RI_ACC[13] ), .B(\pk_rwrit_h[68] ) );
    snl_ao023x1 \REGF/pbmemff11/U883  ( .Z(\REGF/pbmemff11/RO_STAT5BP[3] ), 
        .A(\REGF/pbmemff11/n5136 ), .B(\REGF/pbmemff11/n5137 ), .C(
        \pk_stat_h[18] ), .D(\REGF/RI_STAT[3] ), .E(\REGF/pbmemff11/n5138 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[22]  ( .Q(\pk_indy_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDY389[22] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U913  ( .ZN(\REGF/pbmemff11/n5121 ), .A(PDLIN
        [17]) );
    snl_and02x1 \REGF/pbmemff11/U693  ( .Z(\REGF/pbmemff11/RO_ACC147[30] ), 
        .A(\REGF/RI_ACC[30] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U703  ( .ZN(\REGF/pbmemff11/RO_INDW309[8] ), 
        .A(\REGF/pbmemff11/n5112 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U808  ( .ZN(\REGF/pbmemff11/RO_INDY389[21] ), 
        .A(\REGF/pbmemff11/n5125 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U841  ( .ZN(\REGF/pbmemff11/RO_INDX349[22] ), 
        .A(\REGF/pbmemff11/n5126 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U724  ( .ZN(\REGF/pbmemff11/RO_INDW309[29] ), 
        .A(\REGF/pbmemff11/n5133 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U788  ( .ZN(\REGF/pbmemff11/RO_INDY389[1] ), 
        .A(\REGF/pbmemff11/n5105 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U866  ( .ZN(\REGF/pbmemff11/RO_INDZ429[15] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5119 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[21]  ( .Q(\REGF/RO_EACC[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_EACC187[21] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[12]  ( .Q(\REGF/RO_EACC[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[12] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[31]  ( .Q(\REGF/pk_indw_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDW309[31] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[28]  ( .Q(\REGF/pk_indw_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDW309[28] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[10]  ( .Q(\pk_indz_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[10] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U636  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[1] ), 
        .A(\REGF/RI_DPR[1] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U643  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[8] ), 
        .A(\REGF/RI_DPR[8] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U681  ( .Z(\REGF/pbmemff11/RO_ACC147[18] ), 
        .A(\REGF/RI_ACC[18] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U853  ( .ZN(\REGF/pbmemff11/RO_INDZ429[2] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5106 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[23]  ( .Q(\pk_indz_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[23] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[8]  ( .Q(\pk_indz_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[8] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_DPR28B_reg[25]  ( .Q(\pk_dpr_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[25] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[16]  ( .Q(\pk_dpr_h[16] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[16] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U711  ( .ZN(\REGF/pbmemff11/RO_INDW309[16] ), 
        .A(\REGF/pbmemff11/n5120 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_and02x1 \REGF/pbmemff11/U736  ( .Z(\REGF/pbmemff11/RO_EACC187[9] ), 
        .A(\pk_rwrit_h[67] ), .B(\REGF/RI_EACC[9] ) );
    snl_and02x1 \REGF/pbmemff11/U758  ( .Z(\REGF/pbmemff11/RO_EACC187[31] ), 
        .A(\REGF/RI_EACC[31] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U874  ( .ZN(\REGF/pbmemff11/RO_INDZ429[23] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5127 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[6]  ( .Q(\pk_spr_h[6] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[6] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[22]  ( .Q(\REGF/RO_ACC[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[22] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[11]  ( .Q(\REGF/RO_ACC[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_ACC147[11] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[5]  ( .Q(\pk_indz_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[5] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[20]  ( .Q(\pk_spr_h[20] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[20] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[13]  ( .Q(\pk_spr_h[13] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[13] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U658  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[23] 
        ), .A(\REGF/RI_DPR[23] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U664  ( .Z(\REGF/pbmemff11/RO_ACC147[1] ), .A(
        \REGF/RI_ACC[1] ), .B(\pk_rwrit_h[68] ) );
    snl_invx05 \REGF/pbmemff11/U891  ( .ZN(\REGF/pbmemff11/n5112 ), .A(PDLIN
        [8]) );
    snl_invx05 \REGF/pbmemff11/U901  ( .ZN(\REGF/pbmemff11/n5132 ), .A(PDLIN
        [28]) );
    snl_nand02x1 \REGF/pbmemff11/U926  ( .ZN(\REGF/pbmemff11/n5143 ), .A(
        \REGF/pbmemff11/n5145 ), .B(\REGF/pbmemff11/n5142 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[25]  ( .Q(\REGF/pk_indw_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDW309[25] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[16]  ( .Q(\pk_indw_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[16] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[18]  ( .Q(\REGF/RO_ACC[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_ACC147[18] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[27]  ( .Q(\REGF/pk_indz_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[27] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[14]  ( .Q(\pk_indz_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[14] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U743  ( .Z(\REGF/pbmemff11/RO_EACC187[16] ), 
        .A(\REGF/RI_EACC[16] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U764  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[5] ), 
        .A(\REGF/RI_SPR[5] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[25]  ( .Q(\REGF/RO_EACC[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_EACC187[25] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U801  ( .ZN(\REGF/pbmemff11/RO_INDY389[14] ), 
        .A(\REGF/pbmemff11/n5118 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U826  ( .ZN(\REGF/pbmemff11/RO_INDX349[7] ), 
        .A(\REGF/pbmemff11/n5111 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[16]  ( .Q(\REGF/RO_EACC[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[16] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U848  ( .ZN(\REGF/pbmemff11/RO_INDX349[29] ), 
        .A(\REGF/pbmemff11/n5133 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_invx2 \REGF/pbmemff11/U612  ( .ZN(\REGF/pbmemff11/n5092 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_ffqsnx1 \REGF/pbmemff11/RO_STAT5B_reg[2]  ( .Q(\REGF/pk_stat_h[16] ), 
        .D(pk_ciffh), .SN(\REGF/pbmemff11/n5090 ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff11/U613  ( .ZN(\REGF/pbmemff11/n5086 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_invx1 \REGF/pbmemff11/U626  ( .ZN(\REGF/pbmemff11/n5097 ), .A(
        \REGF/pbmemff11/n5096 ) );
    snl_nand12x1 \REGF/pbmemff11/U648  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[13] 
        ), .A(\REGF/RI_DPR[13] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U653  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[18] 
        ), .A(\REGF/RI_DPR[18] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U674  ( .Z(\REGF/pbmemff11/RO_ACC147[11] ), 
        .A(\REGF/RI_ACC[11] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U691  ( .Z(\REGF/pbmemff11/RO_ACC147[28] ), 
        .A(\REGF/RI_ACC[28] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U701  ( .ZN(\REGF/pbmemff11/RO_INDW309[6] ), 
        .A(\REGF/pbmemff11/n5110 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U726  ( .ZN(\REGF/pbmemff11/RO_INDW309[31] ), 
        .A(\REGF/pbmemff11/n5135 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nand12x1 \REGF/pbmemff11/U781  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[22] 
        ), .A(\REGF/RI_SPR[22] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[26]  ( .Q(\REGF/pk_indy_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDY389[26] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[15]  ( .Q(\pk_indy_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[15] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_DPR28B_reg[24]  ( .Q(\pk_dpr_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[24] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[17]  ( .Q(\pk_dpr_h[17] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[17] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U843  ( .ZN(\REGF/pbmemff11/RO_INDX349[24] ), 
        .A(\REGF/pbmemff11/n5128 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U864  ( .ZN(\REGF/pbmemff11/RO_INDZ429[13] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5117 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[7]  ( .Q(\pk_spr_h[7] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[7] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U748  ( .Z(\REGF/pbmemff11/RO_EACC187[21] ), 
        .A(\REGF/RI_EACC[21] ), .B(\pk_rwrit_h[67] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[23]  ( .Q(\REGF/RO_ACC[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[23] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[10]  ( .Q(\REGF/RO_ACC[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[10] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[4]  ( .Q(\pk_indz_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[4] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[21]  ( .Q(\pk_spr_h[21] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[21] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[12]  ( .Q(\pk_spr_h[12] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[12] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[24]  ( .Q(\REGF/pk_indw_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDW309[24] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[17]  ( .Q(\pk_indw_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDW309[17] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U881  ( .ZN(\REGF/pbmemff11/RO_INDZ429[30] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5134 ) );
    snl_invx05 \REGF/pbmemff11/U911  ( .ZN(\REGF/pbmemff11/n5123 ), .A(PDLIN
        [19]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[26]  ( .Q(\REGF/pk_indz_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[26] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[15]  ( .Q(\pk_indz_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[15] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U753  ( .Z(\REGF/pbmemff11/RO_EACC187[26] ), 
        .A(\REGF/RI_EACC[26] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U811  ( .ZN(\REGF/pbmemff11/RO_INDY389[24] ), 
        .A(\REGF/pbmemff11/n5128 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[19]  ( .Q(\REGF/RO_ACC[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[19] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_nand12x1 \REGF/pbmemff11/U774  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[15] 
        ), .A(\REGF/RI_SPR[15] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U791  ( .ZN(\REGF/pbmemff11/RO_INDY389[4] ), 
        .A(\REGF/pbmemff11/n5108 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U836  ( .ZN(\REGF/pbmemff11/RO_INDX349[17] ), 
        .A(\REGF/pbmemff11/n5121 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[24]  ( .Q(\REGF/RO_EACC[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[24] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U858  ( .ZN(\REGF/pbmemff11/RO_INDZ429[7] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5111 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[17]  ( .Q(\REGF/RO_EACC[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_EACC187[17] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[14]  ( .Q(\pk_indy_h[14] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDY389[14] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[27]  ( .Q(\REGF/pk_indy_h[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDY389[27] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_invx2 \REGF/pbmemff11/U614  ( .ZN(\REGF/pbmemff11/n5088 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_invx1 \REGF/pbmemff11/U628  ( .ZN(\REGF/pbmemff11/n5099 ), .A(
        \REGF/pbmemff11/n5098 ) );
    snl_nand02x1 \REGF/pbmemff11/U634  ( .ZN(\REGF/pbmemff11/n_4044 ), .A(
        \REGF/pbmemff11/n5102 ), .B(\REGF/pbmemff11/n5643 ) );
    snl_and02x1 \REGF/pbmemff11/U783  ( .Z(\REGF/pbmemff11/RO_SPR28B268[24] ), 
        .A(\REGF/RI_SPR[24] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[30]  ( .Q(\REGF/RO_EACC[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[30] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[20]  ( .Q(\pk_indw_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[20] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[29]  ( .Q(\REGF/RO_EACC[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_EACC187[29] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[13]  ( .Q(\pk_indw_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDW309[13] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U641  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[6] ), 
        .A(\REGF/RI_DPR[6] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U666  ( .Z(\REGF/pbmemff11/RO_ACC147[3] ), .A(
        \REGF/RI_ACC[3] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U698  ( .ZN(\REGF/pbmemff11/RO_INDW309[3] ), 
        .A(\REGF/pbmemff11/n5107 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U708  ( .ZN(\REGF/pbmemff11/RO_INDW309[13] ), 
        .A(\REGF/pbmemff11/n5117 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_and02x1 \REGF/pbmemff11/U741  ( .Z(\REGF/pbmemff11/RO_EACC187[14] ), 
        .A(\REGF/RI_EACC[14] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U803  ( .ZN(\REGF/pbmemff11/RO_INDY389[16] ), 
        .A(\REGF/pbmemff11/n5120 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[27]  ( .Q(\REGF/RO_ACC[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_ACC147[27] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[14]  ( .Q(\REGF/RO_ACC[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_ACC147[14] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[18]  ( .Q(\pk_indz_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[18] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[0]  ( .Q(\pk_indz_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[0] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_SPR28B_reg[25]  ( .Q(\pk_spr_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[25] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[16]  ( .Q(\pk_spr_h[16] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[16] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U766  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[7] ), 
        .A(\REGF/RI_SPR[7] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[19]  ( .Q(\pk_indy_h[19] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[19] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U824  ( .ZN(\REGF/pbmemff11/RO_INDX349[5] ), 
        .A(\REGF/pbmemff11/n5109 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[3]  ( .Q(\pk_spr_h[3] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[3] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U888  ( .ZN(\REGF/pbmemff11/n5144 ), .A(
        ph_ciwt_h), .B(\pk_rwrit_h[60] ) );
    snl_invx05 \REGF/pbmemff11/U918  ( .ZN(\REGF/pbmemff11/n5116 ), .A(PDLIN
        [12]) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[13]  ( .Q(\pk_dpr_h[13] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[13] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U924  ( .ZN(\REGF/pbmemff11/n5140 ), .A(
        ph_ebaccwt_h) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[20]  ( .Q(\pk_dpr_h[20] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[20] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U683  ( .Z(\REGF/pbmemff11/RO_ACC147[20] ), 
        .A(\REGF/RI_ACC[20] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U734  ( .Z(\REGF/pbmemff11/RO_EACC187[7] ), 
        .A(\REGF/RI_EACC[7] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U818  ( .ZN(\REGF/pbmemff11/RO_INDY389[31] ), 
        .A(\REGF/pbmemff11/n5135 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_invx05 \REGF/pbmemff11/U893  ( .ZN(\REGF/pbmemff11/n5110 ), .A(PDLIN
        [6]) );
    snl_invx05 \REGF/pbmemff11/U903  ( .ZN(\REGF/pbmemff11/n5130 ), .A(PDLIN
        [26]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[10]  ( .Q(\pk_indy_h[10] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDY389[10] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[23]  ( .Q(\pk_indy_h[23] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[23] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[20]  ( .Q(\REGF/RO_EACC[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[20] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U851  ( .ZN(\REGF/pbmemff11/RO_INDZ429[0] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5104 ) );
    snl_nor02x1 \REGF/pbmemff11/U876  ( .ZN(\REGF/pbmemff11/RO_INDZ429[25] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5129 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[13]  ( .Q(\REGF/RO_EACC[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_EACC187[13] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[30]  ( .Q(\REGF/pk_indw_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDW309[30] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[29]  ( .Q(\REGF/pk_indw_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDW309[29] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U684  ( .Z(\REGF/pbmemff11/RO_ACC147[21] ), 
        .A(\REGF/RI_ACC[21] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U713  ( .ZN(\REGF/pbmemff11/RO_INDW309[18] ), 
        .A(\REGF/pbmemff11/n5122 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U714  ( .ZN(\REGF/pbmemff11/RO_INDW309[19] ), 
        .A(\REGF/pbmemff11/n5123 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U798  ( .ZN(\REGF/pbmemff11/RO_INDY389[11] ), 
        .A(\REGF/pbmemff11/n5115 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[11]  ( .Q(\pk_indz_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[11] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[9]  ( .Q(\pk_indz_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[9] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[22]  ( .Q(\pk_indz_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[22] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U733  ( .Z(\REGF/pbmemff11/RO_EACC187[6] ), 
        .A(\REGF/RI_EACC[6] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U856  ( .ZN(\REGF/pbmemff11/RO_INDZ429[5] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5109 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[22]  ( .Q(\REGF/RO_EACC[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_EACC187[22] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[18]  ( .Q(\pk_indw_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDW309[18] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U871  ( .ZN(\REGF/pbmemff11/RO_INDZ429[20] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5124 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[11]  ( .Q(\REGF/RO_EACC[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_EACC187[11] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[20]  ( .Q(\pk_indz_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[20] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[13]  ( .Q(\pk_indz_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[13] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_nand02x1 \REGF/pbmemff11/U633  ( .ZN(\REGF/pbmemff11/n_3464 ), .A(
        \REGF/pbmemff11/n5101 ), .B(\REGF/pbmemff11/n5643 ) );
    snl_nand12x1 \REGF/pbmemff11/U646  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[11] 
        ), .A(\REGF/RI_DPR[11] ), .B(\pk_rwrit_h[66] ) );
    snl_invx05 \REGF/pbmemff11/U894  ( .ZN(\REGF/pbmemff11/n5109 ), .A(PDLIN
        [5]) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[8]  ( .Q(\pk_spr_h[8] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[8] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_invx05 \REGF/pbmemff11/U904  ( .ZN(\REGF/pbmemff11/n5129 ), .A(PDLIN
        [25]) );
    snl_and02x1 \REGF/pbmemff11/U661  ( .Z(\REGF/pbmemff11/RO_DPR28B227[26] ), 
        .A(\REGF/RI_DPR[26] ), .B(\pk_rwrit_h[66] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[12]  ( .Q(\pk_indy_h[12] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[12] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U746  ( .Z(\REGF/pbmemff11/RO_EACC187[19] ), 
        .A(\REGF/RI_EACC[19] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U761  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[2] ), 
        .A(\REGF/RI_SPR[2] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U823  ( .ZN(\REGF/pbmemff11/RO_INDX349[4] ), 
        .A(\REGF/pbmemff11/n5108 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U838  ( .ZN(\REGF/pbmemff11/RO_INDX349[19] ), 
        .A(\REGF/pbmemff11/n5123 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_invx05 \REGF/pbmemff11/U923  ( .ZN(\REGF/pbmemff11/n5137 ), .A(
        ph_ltwt_h) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[21]  ( .Q(\pk_indy_h[21] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[21] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[31]  ( .Q(\REGF/pk_indy_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDY389[31] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[28]  ( .Q(\REGF/pk_indy_h[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDY389[28] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[18]  ( .Q(\pk_dpr_h[18] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[18] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U804  ( .ZN(\REGF/pbmemff11/RO_INDY389[17] ), 
        .A(\REGF/pbmemff11/n5121 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[22]  ( .Q(\pk_dpr_h[22] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[22] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[11]  ( .Q(\pk_dpr_h[11] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[11] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[1]  ( .Q(\pk_spr_h[1] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[1] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U784  ( .Z(\REGF/pbmemff11/RO_SPR28B268[25] ), 
        .A(\REGF/RI_SPR[25] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[18]  ( .Q(\REGF/RO_EACC[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_EACC187[18] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[22]  ( .Q(\pk_indw_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDW309[22] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_invx2 \REGF/pbmemff11/U615  ( .ZN(\REGF/pbmemff11/n5087 ), .A(
        \REGF/pbmemff11/n5089 ) );
    snl_nand12x8 \REGF/pbmemff11/U621  ( .ZN(\REGF/pbmemff11/n_452 ), .A(
        \pk_rwrit_h[68] ), .B(\REGF/pbmemff11/n5643 ) );
    snl_and02x1 \REGF/pbmemff11/U728  ( .Z(\REGF/pbmemff11/RO_EACC187[1] ), 
        .A(\REGF/RI_EACC[1] ), .B(\pk_rwrit_h[67] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[11]  ( .Q(\pk_indw_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[11] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[30]  ( .Q(\REGF/pk_indz_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[30] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[29]  ( .Q(\REGF/pk_indz_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[29] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U878  ( .ZN(\REGF/pbmemff11/RO_INDZ429[27] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5131 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[25]  ( .Q(\REGF/RO_ACC[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_ACC147[25] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[16]  ( .Q(\REGF/RO_ACC[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_ACC147[16] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[2]  ( .Q(\pk_indz_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[2] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_SPR28B_reg[27]  ( .Q(\pk_spr_h[31] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[27] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[14]  ( .Q(\pk_spr_h[14] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[14] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_invx1 \REGF/pbmemff11/U632  ( .ZN(\REGF/pbmemff11/n5103 ), .A(
        \pk_rwrit_h[61] ) );
    snl_nand12x1 \REGF/pbmemff11/U654  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[19] 
        ), .A(\REGF/RI_DPR[19] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U668  ( .Z(\REGF/pbmemff11/RO_ACC147[5] ), .A(
        \REGF/RI_ACC[5] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U796  ( .ZN(\REGF/pbmemff11/RO_INDY389[9] ), 
        .A(\REGF/pbmemff11/n5113 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[25]  ( .Q(\REGF/pk_indy_h[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDY389[25] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[16]  ( .Q(\pk_indy_h[16] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[16] ), .SE(\REGF/pbmemff11/n5094 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[17]  ( .Q(\pk_indz_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[17] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U754  ( .Z(\REGF/pbmemff11/RO_EACC187[27] ), 
        .A(\REGF/RI_EACC[27] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U773  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[14] 
        ), .A(\REGF/RI_SPR[14] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U831  ( .ZN(\REGF/pbmemff11/RO_INDX349[12] ), 
        .A(\REGF/pbmemff11/n5116 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[31]  ( .Q(pk_sign_h), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_ACC147[31] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[24]  ( .Q(\REGF/pk_indz_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[24] ), .SE(\REGF/pbmemff11/n5099 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[19]  ( .Q(\pk_spr_h[19] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[19] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[28]  ( .Q(\REGF/RO_ACC[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_ACC147[28] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[26]  ( .Q(\REGF/RO_EACC[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[26] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U768  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[9] ), 
        .A(\REGF/RI_SPR[9] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U816  ( .ZN(\REGF/pbmemff11/RO_INDY389[29] ), 
        .A(\REGF/pbmemff11/n5133 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[15]  ( .Q(\REGF/RO_EACC[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_EACC187[15] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[21]  ( .Q(\REGF/RO_ACC[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_ACC147[21] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[12]  ( .Q(\REGF/RO_ACC[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_ACC147[12] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK
        ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[23]  ( .Q(\pk_spr_h[23] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[23] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDZ_reg[6]  ( .Q(\pk_indz_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDZ429[6] ), .SE(\REGF/pbmemff11/n5099 ), .CP(SCLK
        ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[10]  ( .Q(\pk_spr_h[10] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[10] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_ao023x1 \REGF/pbmemff11/U886  ( .Z(pk_bacch), .A(
        \REGF/pbmemff11/n5136 ), .B(\REGF/pbmemff11/n5142 ), .C(\pk_stat_h[0] 
        ), .D(\REGF/RI_STAT[0] ), .E(\REGF/pbmemff11/n5143 ) );
    snl_invx05 \REGF/pbmemff11/U916  ( .ZN(\REGF/pbmemff11/n5118 ), .A(PDLIN
        [14]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[26]  ( .Q(\REGF/pk_indw_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDW309[26] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[15]  ( .Q(\pk_indw_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDW309[15] ), .SE(\REGF/pbmemff11/n5097 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U673  ( .Z(\REGF/pbmemff11/RO_ACC147[10] ), 
        .A(\REGF/RI_ACC[10] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U696  ( .ZN(\REGF/pbmemff11/RO_INDW309[1] ), 
        .A(\REGF/pbmemff11/n5105 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_DPR28B_reg[26]  ( .Q(\pk_dpr_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[26] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[15]  ( .Q(\pk_dpr_h[15] ), 
        .D(1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[15] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U706  ( .ZN(\REGF/pbmemff11/RO_INDW309[11] ), 
        .A(\REGF/pbmemff11/n5115 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U721  ( .ZN(\REGF/pbmemff11/RO_INDW309[26] ), 
        .A(\REGF/pbmemff11/n5130 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U844  ( .ZN(\REGF/pbmemff11/RO_INDX349[25] ), 
        .A(\REGF/pbmemff11/n5129 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_SPR28B_reg[5]  ( .Q(\pk_spr_h[5] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_SPR28B268[5] ), .SE(\REGF/pbmemff11/n_2192 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U863  ( .ZN(\REGF/pbmemff11/RO_INDZ429[12] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5116 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[2]  ( .Q(\REGF/RO_EACC[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_EACC187[2] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[9]  ( .Q(\pk_dpr_h[9] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[9] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_invx1 \REGF/pbmemff11/U629  ( .ZN(\REGF/pbmemff11/n5101 ), .A(
        \pk_rwrit_h[63] ) );
    snl_nand12x1 \REGF/pbmemff11/U647  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[12] 
        ), .A(\REGF/RI_DPR[12] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U729  ( .Z(\REGF/pbmemff11/RO_EACC187[2] ), 
        .A(\REGF/RI_EACC[2] ), .B(\pk_rwrit_h[67] ) );
    snl_and02x1 \REGF/pbmemff11/U785  ( .Z(\REGF/pbmemff11/RO_SPR28B268[26] ), 
        .A(\REGF/RI_SPR[26] ), .B(\pk_rwrit_h[65] ) );
    snl_and02x1 \REGF/pbmemff11/U747  ( .Z(\REGF/pbmemff11/RO_EACC187[20] ), 
        .A(\REGF/RI_EACC[20] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U760  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[1] ), 
        .A(\REGF/RI_SPR[1] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U822  ( .ZN(\REGF/pbmemff11/RO_INDX349[3] ), 
        .A(\REGF/pbmemff11/n5107 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[0]  ( .Q(\REGF/RO_ACC[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_ACC147[0] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_nor02x1 \REGF/pbmemff11/U805  ( .ZN(\REGF/pbmemff11/RO_INDY389[18] ), 
        .A(\REGF/pbmemff11/n5122 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_invx05 \REGF/pbmemff11/U895  ( .ZN(\REGF/pbmemff11/n5108 ), .A(PDLIN
        [4]) );
    snl_invx05 \REGF/pbmemff11/U905  ( .ZN(\REGF/pbmemff11/n5128 ), .A(PDLIN
        [24]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[9]  ( .Q(\pk_indw_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDW309[9] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_and02x1 \REGF/pbmemff11/U660  ( .Z(\REGF/pbmemff11/RO_DPR28B227[25] ), 
        .A(\REGF/RI_DPR[25] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U685  ( .Z(\REGF/pbmemff11/RO_ACC147[22] ), 
        .A(\REGF/RI_ACC[22] ), .B(\pk_rwrit_h[68] ) );
    snl_nor02x1 \REGF/pbmemff11/U839  ( .ZN(\REGF/pbmemff11/RO_INDX349[20] ), 
        .A(\REGF/pbmemff11/n5124 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_invx05 \REGF/pbmemff11/U922  ( .ZN(\REGF/pbmemff11/n5145 ), .A(
        \pk_rwrit_h[60] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[0]  ( .Q(\pk_indw_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDW309[0] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[5]  ( .Q(\pk_indy_h[5] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDY389[5] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[26]  ( .Q(\REGF/pk_indx_h[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDX349[26] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U715  ( .ZN(\REGF/pbmemff11/RO_INDW309[20] ), 
        .A(\REGF/pbmemff11/n5124 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_and02x1 \REGF/pbmemff11/U732  ( .Z(\REGF/pbmemff11/RO_EACC187[5] ), 
        .A(\REGF/RI_EACC[5] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U857  ( .ZN(\REGF/pbmemff11/RO_INDZ429[6] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5110 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[15]  ( .Q(\pk_indx_h[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[15] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[0]  ( .Q(\pk_dpr_h[0] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[0] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U870  ( .ZN(\REGF/pbmemff11/RO_INDZ429[19] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5123 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[9]  ( .Q(\REGF/RO_ACC[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_ACC147[9] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_nand12x1 \REGF/pbmemff11/U655  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[20] 
        ), .A(\REGF/RI_DPR[20] ), .B(\pk_rwrit_h[66] ) );
    snl_nor02x1 \REGF/pbmemff11/U697  ( .ZN(\REGF/pbmemff11/RO_INDW309[2] ), 
        .A(\REGF/pbmemff11/n5106 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U707  ( .ZN(\REGF/pbmemff11/RO_INDW309[12] ), 
        .A(\REGF/pbmemff11/n5116 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[2]  ( .Q(\pk_indx_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDX349[2] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[8]  ( .Q(\pk_indy_h[8] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDY389[8] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_nor02x1 \REGF/pbmemff11/U720  ( .ZN(\REGF/pbmemff11/RO_INDW309[25] ), 
        .A(\REGF/pbmemff11/n5129 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U845  ( .ZN(\REGF/pbmemff11/RO_INDX349[26] ), 
        .A(\REGF/pbmemff11/n5130 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U862  ( .ZN(\REGF/pbmemff11/RO_INDZ429[11] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5115 ) );
    snl_nand12x1 \REGF/pbmemff11/U769  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[10] 
        ), .A(\REGF/RI_SPR[10] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[4]  ( .Q(\REGF/RO_ACC[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_ACC147[4] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_invx05 \REGF/pbmemff11/U887  ( .ZN(\REGF/pbmemff11/n5643 ), .A(
        \pk_rwrit_h[44] ) );
    snl_invx05 \REGF/pbmemff11/U917  ( .ZN(\REGF/pbmemff11/n5117 ), .A(PDLIN
        [13]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[18]  ( .Q(\pk_indx_h[18] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDX349[18] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U669  ( .Z(\REGF/pbmemff11/RO_ACC147[6] ), .A(
        \REGF/RI_ACC[6] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U672  ( .Z(\REGF/pbmemff11/RO_ACC147[9] ), .A(
        \pk_rwrit_h[68] ), .B(\REGF/RI_ACC[9] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[6]  ( .Q(\REGF/RO_EACC[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_EACC187[6] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[6]  ( .Q(\pk_indx_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDX349[6] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_and02x1 \REGF/pbmemff11/U755  ( .Z(\REGF/pbmemff11/RO_EACC187[28] ), 
        .A(\REGF/RI_EACC[28] ), .B(\pk_rwrit_h[67] ) );
    snl_nand12x1 \REGF/pbmemff11/U772  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[13] 
        ), .A(\REGF/RI_SPR[13] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U830  ( .ZN(\REGF/pbmemff11/RO_INDX349[11] ), 
        .A(\REGF/pbmemff11/n5115 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U817  ( .ZN(\REGF/pbmemff11/RO_INDY389[30] ), 
        .A(\REGF/pbmemff11/n5134 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[22]  ( .Q(\pk_indx_h[22] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[22] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U879  ( .ZN(\REGF/pbmemff11/RO_INDZ429[28] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5132 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[11]  ( .Q(\pk_indx_h[11] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDX349[11] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[4]  ( .Q(\pk_dpr_h[4] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[4] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[1]  ( .Q(\pk_indy_h[1] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[1] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[4]  ( .Q(\pk_indw_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDW309[4] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_nand12x8 \REGF/pbmemff11/U620  ( .ZN(\REGF/pbmemff11/n_2192 ), .A(
        \pk_rwrit_h[65] ), .B(\REGF/pbmemff11/n5643 ) );
    snl_and02x1 \REGF/pbmemff11/U627  ( .Z(\REGF/pbmemff11/n5098 ), .A(
        \REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5643 ) );
    snl_nor02x1 \REGF/pbmemff11/U790  ( .ZN(\REGF/pbmemff11/RO_INDY389[3] ), 
        .A(\REGF/pbmemff11/n5107 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U797  ( .ZN(\REGF/pbmemff11/RO_INDY389[10] ), 
        .A(\REGF/pbmemff11/n5114 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U859  ( .ZN(\REGF/pbmemff11/RO_INDZ429[8] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5112 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[3]  ( .Q(\pk_indy_h[3] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[3] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[6]  ( .Q(\pk_indw_h[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_INDW309[6] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_ffqrnx1 \REGF/pbmemff11/RO_STAT5B_reg[0]  ( .Q(\pk_stat_h[0] ), .D(
        pk_bacch), .RN(\REGF/pbmemff11/n5092 ), .CP(SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U640  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[5] ), 
        .A(\REGF/RI_DPR[5] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U649  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[14] 
        ), .A(\REGF/RI_DPR[14] ), .B(\pk_rwrit_h[66] ) );
    snl_nand12x1 \REGF/pbmemff11/U652  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[17] 
        ), .A(\REGF/RI_DPR[17] ), .B(\pk_rwrit_h[66] ) );
    snl_and02x1 \REGF/pbmemff11/U675  ( .Z(\REGF/pbmemff11/RO_ACC147[12] ), 
        .A(\REGF/RI_ACC[12] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U749  ( .Z(\REGF/pbmemff11/RO_EACC187[22] ), 
        .A(\REGF/RI_EACC[22] ), .B(\pk_rwrit_h[67] ) );
    snl_and02x1 \REGF/pbmemff11/U752  ( .Z(\REGF/pbmemff11/RO_EACC187[25] ), 
        .A(\REGF/RI_EACC[25] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U810  ( .ZN(\REGF/pbmemff11/RO_INDY389[23] ), 
        .A(\REGF/pbmemff11/n5127 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[4]  ( .Q(\pk_indx_h[4] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_INDX349[4] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_nand12x1 \REGF/pbmemff11/U775  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[16] 
        ), .A(\REGF/RI_SPR[16] ), .B(\pk_rwrit_h[65] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[20]  ( .Q(\pk_indx_h[20] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_INDX349[20] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U837  ( .ZN(\REGF/pbmemff11/RO_INDX349[18] ), 
        .A(\REGF/pbmemff11/n5122 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[13]  ( .Q(\pk_indx_h[13] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDX349[13] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[6]  ( .Q(\pk_dpr_h[6] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[6] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[6]  ( .Q(\REGF/RO_ACC[6] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_ACC147[6] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[30]  ( .Q(\REGF/pk_indx_h[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5090 ), .SD(
        \REGF/pbmemff11/RO_INDX349[30] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[29]  ( .Q(\REGF/pk_indx_h[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDX349[29] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[4]  ( .Q(\REGF/RO_EACC[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5088 ), .SD(
        \REGF/pbmemff11/RO_EACC187[4] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_and02x1 \REGF/pbmemff11/U667  ( .Z(\REGF/pbmemff11/RO_ACC147[4] ), .A(
        \REGF/RI_ACC[4] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U682  ( .Z(\REGF/pbmemff11/RO_ACC147[19] ), 
        .A(\REGF/RI_ACC[19] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U690  ( .Z(\REGF/pbmemff11/RO_ACC147[27] ), 
        .A(\REGF/RI_ACC[27] ), .B(\pk_rwrit_h[68] ) );
    snl_and02x1 \REGF/pbmemff11/U727  ( .Z(\REGF/pbmemff11/RO_EACC187[0] ), 
        .A(\REGF/RI_EACC[0] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U880  ( .ZN(\REGF/pbmemff11/RO_INDZ429[29] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5133 ) );
    snl_invx05 \REGF/pbmemff11/U910  ( .ZN(\REGF/pbmemff11/n5105 ), .A(PDLIN
        [1]) );
    snl_nor02x1 \REGF/pbmemff11/U842  ( .ZN(\REGF/pbmemff11/RO_INDX349[23] ), 
        .A(\REGF/pbmemff11/n5127 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U865  ( .ZN(\REGF/pbmemff11/RO_INDZ429[14] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5118 ) );
    snl_nor02x1 \REGF/pbmemff11/U700  ( .ZN(\REGF/pbmemff11/RO_INDW309[5] ), 
        .A(\REGF/pbmemff11/n5109 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U712  ( .ZN(\REGF/pbmemff11/RO_INDW309[17] ), 
        .A(\REGF/pbmemff11/n5121 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_and02x1 \REGF/pbmemff11/U735  ( .Z(\REGF/pbmemff11/RO_EACC187[8] ), 
        .A(\REGF/RI_EACC[8] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U850  ( .ZN(\REGF/pbmemff11/RO_INDX349[31] ), 
        .A(\REGF/pbmemff11/n5135 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U877  ( .ZN(\REGF/pbmemff11/RO_INDZ429[26] ), 
        .A(\REGF/pbmemff11/n5103 ), .B(\REGF/pbmemff11/n5130 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[24]  ( .Q(\REGF/pk_indx_h[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[24] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[17]  ( .Q(\pk_indx_h[17] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[17] ), .SE(\REGF/pbmemff11/n5095 ), .CP(
        SCLK) );
    snl_sffqensnx2 \REGF/pbmemff11/RO_DPR28B_reg[2]  ( .Q(\pk_dpr_h[2] ), .D(
        1'b0), .EN(1'b1), .SN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_DPR28B227[2] ), .SE(\REGF/pbmemff11/n_1556 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U799  ( .ZN(\REGF/pbmemff11/RO_INDY389[12] ), 
        .A(\REGF/pbmemff11/n5116 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[9]  ( .Q(\REGF/RO_EACC[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_EACC187[9] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[0]  ( .Q(\pk_indx_h[0] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[0] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_invx05 \REGF/pbmemff11/U925  ( .ZN(\REGF/pbmemff11/n5142 ), .A(
        ph_baccwt_h) );
    snl_and02x1 \REGF/pbmemff11/U740  ( .Z(\REGF/pbmemff11/RO_EACC187[13] ), 
        .A(\REGF/RI_EACC[13] ), .B(\pk_rwrit_h[67] ) );
    snl_nor02x1 \REGF/pbmemff11/U802  ( .ZN(\REGF/pbmemff11/RO_INDY389[15] ), 
        .A(\REGF/pbmemff11/n5119 ), .B(\REGF/pbmemff11/n5102 ) );
    snl_nor02x1 \REGF/pbmemff11/U819  ( .ZN(\REGF/pbmemff11/RO_INDX349[0] ), 
        .A(\REGF/pbmemff11/n5104 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_invx05 \REGF/pbmemff11/U892  ( .ZN(\REGF/pbmemff11/n5111 ), .A(PDLIN
        [7]) );
    snl_invx05 \REGF/pbmemff11/U902  ( .ZN(\REGF/pbmemff11/n5131 ), .A(PDLIN
        [27]) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDW_reg[2]  ( .Q(\pk_indw_h[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5091 ), .SD(
        \REGF/pbmemff11/RO_INDW309[2] ), .SE(\REGF/pbmemff11/n5097 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDY_reg[7]  ( .Q(\pk_indy_h[7] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5087 ), .SD(
        \REGF/pbmemff11/RO_INDY389[7] ), .SE(\REGF/pbmemff11/n5094 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_STAT5B_reg[4]  ( .Q(\REGF/pk_stat_h[30] 
        ), .D(1'b0), .EN(\REGF/pbmemff11/n5643 ), .RN(\REGF/pbmemff11/n5090 ), 
        .SD(\REGF/RI_STAT[4] ), .SE(\pk_rwrit_h[60] ), .CP(SCLK) );
    snl_nand12x1 \REGF/pbmemff11/U767  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[8] ), 
        .A(\REGF/RI_SPR[8] ), .B(\pk_rwrit_h[65] ) );
    snl_nand12x1 \REGF/pbmemff11/U782  ( .ZN(\REGF/pbmemff11/RO_SPR28B268[23] 
        ), .A(\REGF/RI_SPR[23] ), .B(\pk_rwrit_h[65] ) );
    snl_nor02x1 \REGF/pbmemff11/U825  ( .ZN(\REGF/pbmemff11/RO_INDX349[6] ), 
        .A(\REGF/pbmemff11/n5110 ), .B(\REGF/pbmemff11/n5101 ) );
    snl_nor02x1 \REGF/pbmemff11/U889  ( .ZN(\REGF/pbmemff11/n5136 ), .A(
        \pk_rwrit_h[60] ), .B(\pk_rwrit_h[44] ) );
    snl_invx05 \REGF/pbmemff11/U919  ( .ZN(\REGF/pbmemff11/n5115 ), .A(PDLIN
        [11]) );
    snl_nand12x1 \REGF/pbmemff11/U635  ( .ZN(\REGF/pbmemff11/RO_DPR28B227[0] ), 
        .A(\REGF/RI_DPR[0] ), .B(\pk_rwrit_h[66] ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_EACC_reg[0]  ( .Q(\REGF/RO_EACC[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5093 ), .SD(
        \REGF/pbmemff11/RO_EACC187[0] ), .SE(\REGF/pbmemff11/n_1032 ), .CP(
        SCLK) );
    snl_nor02x1 \REGF/pbmemff11/U699  ( .ZN(\REGF/pbmemff11/RO_INDW309[4] ), 
        .A(\REGF/pbmemff11/n5108 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_nor02x1 \REGF/pbmemff11/U709  ( .ZN(\REGF/pbmemff11/RO_INDW309[14] ), 
        .A(\REGF/pbmemff11/n5118 ), .B(\REGF/pbmemff11/n5100 ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_INDX_reg[9]  ( .Q(\pk_indx_h[9] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5092 ), .SD(
        \REGF/pbmemff11/RO_INDX349[9] ), .SE(\REGF/pbmemff11/n5095 ), .CP(SCLK
        ) );
    snl_sffqenrnx1 \REGF/pbmemff11/RO_ACC_reg[2]  ( .Q(\REGF/RO_ACC[2] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff11/n5086 ), .SD(
        \REGF/pbmemff11/RO_ACC147[2] ), .SE(\REGF/pbmemff11/n_452 ), .CP(SCLK)
         );
    snl_bufx1 \MAIN/ENGIN/U73  ( .Z(\MAIN/ENGIN/n3591 ), .A(\MAIN/n3611 ) );
    snl_nand04x1 \MAIN/ENGIN/U74  ( .ZN(st_exectl), .A(
        \MAIN/ENGIN/a_exectl_st ), .B(\MAIN/ENGIN/b_exectl_st ), .C(
        \MAIN/ENGIN/c_exectl_st ), .D(\MAIN/ENGIN/d_exectl_st ) );
    snl_ao2222x1 \MAIN/ENGIN/U83  ( .Z(\MAIN/decend_en ), .A(
        \MAIN/ENGIN/a_deocenh ), .B(\MAIN/ENGIN/b_dec_stage ), .C(
        \MAIN/ENGIN/d_deocenh ), .D(\MAIN/ENGIN/a_dec_stage ), .E(
        \MAIN/ENGIN/b_deocenh ), .F(\MAIN/ENGIN/c_dec_stage ), .G(
        \MAIN/ENGIN/c_deocenh ), .H(\MAIN/ENGIN/d_dec_stage ) );
    snl_or04x1 \MAIN/ENGIN/U84  ( .Z(\MAIN/st_decctl ), .A(
        \MAIN/ENGIN/b_decctl_st ), .B(\MAIN/ENGIN/d_decctl_st ), .C(
        \MAIN/ENGIN/c_decctl_st ), .D(\MAIN/ENGIN/a_decctl_st ) );
    snl_or02x1 \MAIN/ENGIN/U96  ( .Z(\MAIN/ENGIN/n3594 ), .A(
        \MAIN/b_exec_stage ), .B(\MAIN/d_exec_stage ) );
    snl_ffqnrnx2 \MAIN/ENGIN/exe_temp_reg  ( .QN(\MAIN/ENGIN/n_164 ), .D(
        pk_pexe01_h), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK) );
    snl_nand12x1 \MAIN/ENGIN/U101  ( .ZN(\MAIN/ENGIN/n3603 ), .A(
        \MAIN/ENGIN/a_d2_stage ), .B(\MAIN/ENGIN/n3593 ) );
    snl_or02x1 \MAIN/ENGIN/U91  ( .Z(\MAIN/ENGIN/C_PED4_BR ), .A(
        \MAIN/ENGIN/B_INIT_STAGE ), .B(\MAIN/ENGIN/b_step_end ) );
    snl_aoi022x1 \MAIN/ENGIN/U98  ( .ZN(\MAIN/ENGIN/n3601 ), .A(
        \MAIN/ENGIN/a_cf_stage ), .B(\MAIN/ENGIN/n3602 ), .C(
        \MAIN/ENGIN/c_cf_stage ), .D(\MAIN/ENGIN/n3603 ) );
    snl_sffqenrnx1 \MAIN/ENGIN/a_cf_start2_reg  ( .Q(\MAIN/ENGIN/a_cf_start2 ), 
        .D(1'b0), .EN(\MAIN/ENGIN/n3604 ), .RN(\MAIN/ENGIN/n3591 ), .SD(1'b1), 
        .SE(\MAIN/ENGIN/puls_exec ), .CP(SCLK) );
    snl_nand04x0 \MAIN/ENGIN/U75  ( .ZN(\MAIN/st_swctl ), .A(
        \MAIN/ENGIN/a_swctl_st ), .B(\MAIN/ENGIN/b_swctl_st ), .C(
        \MAIN/ENGIN/c_swctl_st ), .D(\MAIN/ENGIN/d_swctl_st ) );
    snl_or02x1 \MAIN/ENGIN/U82  ( .Z(\MAIN/ENGIN/A_PED4_BR ), .A(
        \MAIN/ENGIN/D_INIT_STAGE ), .B(\MAIN/ENGIN/d_step_end ) );
    snl_invx05 \MAIN/ENGIN/U99  ( .ZN(\MAIN/ENGIN/n3592 ), .A(
        \MAIN/c_exec_stage ) );
    snl_aoi013x0 \MAIN/ENGIN/U90  ( .ZN(cf_wait), .A(\MAIN/ENGIN/n3599 ), .B(
        \MAIN/ENGIN/n3600 ), .C(\MAIN/ENGIN/n3601 ), .D(\MAIN/st_swctl ) );
    snl_or04x1 \MAIN/ENGIN/U85  ( .Z(st_cfctl), .A(\MAIN/ENGIN/a_cfctl_st ), 
        .B(\MAIN/ENGIN/b_cfctl_st ), .C(\MAIN/ENGIN/c_cfctl_st ), .D(
        \MAIN/ENGIN/d_cfctl_st ) );
    snl_nor02x1 \MAIN/ENGIN/U97  ( .ZN(\MAIN/ENGIN/n3597 ), .A(
        \MAIN/c_exec_stage ), .B(\MAIN/a_exec_stage ) );
    snl_invx05 \MAIN/ENGIN/U100  ( .ZN(\MAIN/ENGIN/n3593 ), .A(
        \MAIN/a_exec_stage ) );
    snl_nor02x1 \MAIN/ENGIN/U95  ( .ZN(\MAIN/ENGIN/n3598 ), .A(
        \MAIN/b_exec_stage ), .B(\MAIN/d_exec_stage ) );
    snl_ffqrnx1 \MAIN/ENGIN/WP_PC_reg  ( .Q(\MAIN/WP_PC ), .D(\pk_rwrit_h[59] 
        ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK) );
    snl_ao122x1 \MAIN/ENGIN/U79  ( .Z(\MAIN/ph_rdwr2selh ), .A(
        \MAIN/ENGIN/n3592 ), .B(\MAIN/ENGIN/d_dec_stage ), .C(
        \MAIN/ENGIN/n3593 ), .D(\MAIN/ENGIN/b_dec_stage ), .E(
        \MAIN/ENGIN/n3594 ) );
    snl_oai122x0 \MAIN/ENGIN/U80  ( .ZN(\MAIN/ph_rdwr1selh ), .A(
        \MAIN/b_exec_stage ), .B(\MAIN/ENGIN/n3595 ), .C(\MAIN/d_exec_stage ), 
        .D(\MAIN/ENGIN/n3596 ), .E(\MAIN/ENGIN/n3597 ) );
    snl_or02x1 \MAIN/ENGIN/U87  ( .Z(\MAIN/ENGIN/cf_start ), .A(
        \MAIN/ENGIN/a_cf_start2 ), .B(\MAIN/ENGIN/d_decctl_st ) );
    snl_nand12x1 \MAIN/ENGIN/U102  ( .ZN(\MAIN/ENGIN/n3602 ), .A(
        \MAIN/ENGIN/c_d2_stage ), .B(\MAIN/ENGIN/n3592 ) );
    snl_invx05 \MAIN/ENGIN/U76  ( .ZN(\MAIN/ENGIN/n3607 ), .A(
        \MAIN/ENGIN/dec_st2_rst ) );
    snl_invx05 \MAIN/ENGIN/U77  ( .ZN(\MAIN/ENGIN/n3604 ), .A(
        \MAIN/ENGIN/cf_st2_rst ) );
    snl_and02x1 \MAIN/ENGIN/U89  ( .Z(\MAIN/ENGIN/puls_exec ), .A(pk_pexe01_h), 
        .B(\MAIN/ENGIN/n_164 ) );
    snl_or02x1 \MAIN/ENGIN/U92  ( .Z(\MAIN/ENGIN/dec_start ), .A(
        \MAIN/ENGIN/a_dec_start2 ), .B(\MAIN/ENGIN/a_dec_start ) );
    snl_or02x1 \MAIN/ENGIN/U81  ( .Z(\MAIN/ENGIN/B_PED4_BR ), .A(
        \MAIN/ENGIN/A_INIT_STAGE ), .B(\MAIN/ENGIN/a_step_end ) );
    snl_sffqenrnx1 \MAIN/ENGIN/a_dec_start2_reg  ( .Q(
        \MAIN/ENGIN/a_dec_start2 ), .D(1'b0), .EN(\MAIN/ENGIN/n3607 ), .RN(
        \MAIN/ENGIN/n3591 ), .SD(1'b1), .SE(\MAIN/ENGIN/puls_exec ), .CP(SCLK)
         );
    snl_oai012x1 \MAIN/ENGIN/U104  ( .ZN(\MAIN/ENGIN/n3599 ), .A(
        \MAIN/ENGIN/d_d2_stage ), .B(\MAIN/d_exec_stage ), .C(
        \MAIN/ENGIN/b_cf_stage ) );
    snl_or02x1 \MAIN/ENGIN/U88  ( .Z(\MAIN/ENGIN/D_PED4_BR ), .A(
        \MAIN/ENGIN/C_INIT_STAGE ), .B(\MAIN/ENGIN/c_step_end ) );
    snl_invx05 \MAIN/ENGIN/U93  ( .ZN(\MAIN/ENGIN/n3595 ), .A(
        \MAIN/ENGIN/c_dec_stage ) );
    snl_or04x1 \MAIN/ENGIN/U78  ( .Z(ph_cperr_h), .A(\MAIN/ENGIN/status_wr2 ), 
        .B(\MAIN/ENGIN/status_wr3 ), .C(\MAIN/ENGIN/status_wr4 ), .D(
        \MAIN/ENGIN/status_wr1 ) );
    snl_nand14x0 \MAIN/ENGIN/U86  ( .ZN(ph_rgfile_h), .A(st_exectl), .B(
        \MAIN/ENGIN/n3592 ), .C(\MAIN/ENGIN/n3593 ), .D(\MAIN/ENGIN/n3598 ) );
    snl_invx05 \MAIN/ENGIN/U94  ( .ZN(\MAIN/ENGIN/n3596 ), .A(
        \MAIN/ENGIN/a_dec_stage ) );
    snl_oai012x1 \MAIN/ENGIN/U103  ( .ZN(\MAIN/ENGIN/n3600 ), .A(
        \MAIN/ENGIN/b_d2_stage ), .B(\MAIN/b_exec_stage ), .C(
        \MAIN/ENGIN/d_cf_stage ) );
    snl_invx2 \REGF/pbmemff51/U840  ( .ZN(\REGF/pbmemff51/n4474 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[1]  ( .Q(\pk_s0ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[8]  ( .Q(\pk_s0ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[14]  ( .Q(\pk_s1ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[9]  ( .Q(\pk_s2ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[0]  ( .Q(\pk_s2ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[12]  ( .Q(\pk_s3ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[12]  ( .Q(\pk_s7ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[18]  ( .Q(
        \REGF/pk_scba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[14]  ( .Q(\pk_s5ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[8]  ( .Q(\pk_s9ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[4]  ( .Q(\pk_sbba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[6]  ( .Q(\pk_s7ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[1]  ( .Q(\pk_s9ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[14]  ( .Q(\pk_s8ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[17]  ( .Q(\pk_saba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[3]  ( .Q(\pk_seba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[4]  ( .Q(\pk_s2ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[7]  ( .Q(\pk_s5ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[11]  ( .Q(\pk_scba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[17]  ( .Q(\pk_seba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[10]  ( .Q(\pk_s5ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff51/U837  ( .ZN(\REGF/pbmemff51/n4476 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_invx2 \REGF/pbmemff51/U838  ( .ZN(\REGF/pbmemff51/n4470 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_invx2 \REGF/pbmemff51/U841  ( .ZN(\REGF/pbmemff51/n4472 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[17]  ( .Q(\pk_s0ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[7]  ( .Q(\pk_s0ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[5]  ( .Q(\pk_s0ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[16]  ( .Q(\pk_s3ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[0]  ( .Q(\pk_sbba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[16]  ( .Q(\pk_s7ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[10]  ( .Q(\pk_s1ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[8]  ( .Q(\pk_s5ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[3]  ( .Q(\pk_s5ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[1]  ( .Q(\pk_s5ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[2]  ( .Q(\pk_s7ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[10]  ( .Q(\pk_s8ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[5]  ( .Q(\pk_s9ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[15]  ( .Q(\pk_scba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[13]  ( .Q(\pk_seba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[7]  ( .Q(\pk_seba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[13]  ( .Q(\pk_saba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[9]  ( .Q(\pk_sbba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[0]  ( .Q(\pk_s7ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[12]  ( .Q(\pk_s8ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[7]  ( .Q(\pk_s9ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[11]  ( .Q(\pk_saba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[14]  ( .Q(\pk_s7ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[17]  ( .Q(\pk_scba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[11]  ( .Q(\pk_seba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[5]  ( .Q(\pk_seba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[3]  ( .Q(\pk_s0ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[12]  ( .Q(\pk_s1ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[18]  ( .Q(
        \REGF/pk_seba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[6]  ( .Q(\pk_s2ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[12]  ( .Q(\pk_s5ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[18]  ( .Q(
        \REGF/pk_saba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[2]  ( .Q(\pk_s2ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[14]  ( .Q(\pk_s3ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[9]  ( .Q(\pk_s7ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[10]  ( .Q(\pk_s3ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[5]  ( .Q(\pk_s5ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[2]  ( .Q(\pk_sbba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[13]  ( .Q(\pk_scba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[15]  ( .Q(\pk_seba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[1]  ( .Q(\pk_seba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[4]  ( .Q(\pk_s7ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[16]  ( .Q(\pk_s8ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[3]  ( .Q(\pk_s9ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[15]  ( .Q(\pk_saba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[6]  ( .Q(\pk_sbba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[16]  ( .Q(\pk_s5ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[16]  ( .Q(\pk_s1ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[6]  ( .Q(\pk_s1ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[18]  ( .Q(
        \REGF/pk_s2ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[10]  ( .Q(\pk_s7ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[8]  ( .Q(\pk_seba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[3]  ( .Q(\pk_scba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[12]  ( .Q(\pk_sfba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[7]  ( .Q(\pk_s3ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[8]  ( .Q(\pk_s6ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[17]  ( .Q(\pk_s9ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[9]  ( .Q(\pk_s4ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[14]  ( .Q(\pk_sdba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[18]  ( .Q(
        \REGF/pk_s6ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[12]  ( .Q(\pk_sbba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[2]  ( .Q(\pk_saba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[13]  ( .Q(\pk_s0ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[2]  ( .Q(\pk_s1ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[11]  ( .Q(\pk_s2ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[0]  ( .Q(\pk_s4ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[11]  ( .Q(\pk_s6ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[4]  ( .Q(\pk_sdba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[17]  ( .Q(\pk_s4ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[1]  ( .Q(\pk_s6ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[6]  ( .Q(\pk_s8ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[5]  ( .Q(\pk_sfba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[6]  ( .Q(\pk_saba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[16]  ( .Q(\pk_sbba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[10]  ( .Q(\pk_sdba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[9]  ( .Q(\pk_sdba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[15]  ( .Q(\pk_s2ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[3]  ( .Q(\pk_s3ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[13]  ( .Q(\pk_s4ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[13]  ( .Q(\pk_s9ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[7]  ( .Q(\pk_scba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[16]  ( .Q(\pk_sfba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[8]  ( .Q(\pk_sfba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[5]  ( .Q(\pk_s6ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[2]  ( .Q(\pk_s8ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[1]  ( .Q(\pk_sfba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[4]  ( .Q(\pk_s4ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[15]  ( .Q(\pk_s6ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[11]  ( .Q(\pk_s0ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[9]  ( .Q(\pk_s1ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[6]  ( .Q(\pk_s4ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[17]  ( .Q(\pk_s6ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[0]  ( .Q(\pk_sdba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[17]  ( .Q(\pk_s2ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[8]  ( .Q(\pk_s3ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[11]  ( .Q(\pk_s4ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[2]  ( .Q(\pk_sdba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[3]  ( .Q(\pk_sfba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[18]  ( .Q(
        \REGF/pk_s9ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[0]  ( .Q(\pk_s8ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[1]  ( .Q(\pk_s3ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[7]  ( .Q(\pk_s6ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[18]  ( .Q(
        \REGF/pk_s4ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[9]  ( .Q(\pk_s8ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[11]  ( .Q(\pk_s9ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[5]  ( .Q(\pk_scba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[14]  ( .Q(\pk_sfba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff51/U843  ( .ZN(\REGF/pbmemff51/n4475 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[18]  ( .Q(
        \REGF/pk_s0ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[4]  ( .Q(\pk_saba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[14]  ( .Q(\pk_sbba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[12]  ( .Q(\pk_sdba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[15]  ( .Q(\pk_s0ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[0]  ( .Q(\pk_s1ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[13]  ( .Q(\pk_s2ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[3]  ( .Q(\pk_s6ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[15]  ( .Q(\pk_s4ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[4]  ( .Q(\pk_s8ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[8]  ( .Q(\pk_scba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[7]  ( .Q(\pk_sfba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[4]  ( .Q(\pk_s1ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[2]  ( .Q(\pk_s4ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[13]  ( .Q(\pk_s6ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[9]  ( .Q(\pk_saba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[6]  ( .Q(\pk_sdba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[0]  ( .Q(\pk_saba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[10]  ( .Q(\pk_sbba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[16]  ( .Q(\pk_sdba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[1]  ( .Q(\pk_scba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[10]  ( .Q(\pk_sfba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[12]  ( .Q(\pk_s2ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[5]  ( .Q(\pk_s3ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[15]  ( .Q(\pk_s9ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[9]  ( .Q(\pk_scba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[14]  ( .Q(\pk_s4ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[2]  ( .Q(\pk_s6ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[18]  ( .Q(
        \REGF/pk_sfba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[5]  ( .Q(\pk_s8ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[6]  ( .Q(\pk_sfba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[14]  ( .Q(\pk_s0ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[10]  ( .Q(\pk_s0ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[5]  ( .Q(\pk_s1ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[3]  ( .Q(\pk_s4ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[12]  ( .Q(\pk_s6ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[7]  ( .Q(\pk_sdba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[18]  ( .Q(
        \REGF/pk_sbba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[8]  ( .Q(\pk_saba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[17]  ( .Q(\pk_sdba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[4]  ( .Q(\pk_s3ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[1]  ( .Q(\pk_saba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[11]  ( .Q(\pk_sbba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[0]  ( .Q(\pk_scba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[11]  ( .Q(\pk_sfba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[7]  ( .Q(\pk_s4ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[16]  ( .Q(\pk_s6ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[14]  ( .Q(\pk_s9ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[8]  ( .Q(\pk_s1ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[3]  ( .Q(\pk_sdba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[3]  ( .Q(\pk_s1ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[1]  ( .Q(\pk_s1ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[16]  ( .Q(\pk_s2ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[9]  ( .Q(\pk_s3ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[1]  ( .Q(\pk_s8ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[10]  ( .Q(\pk_s4ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[2]  ( .Q(\pk_sfba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[6]  ( .Q(\pk_s6ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[0]  ( .Q(\pk_s3ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[8]  ( .Q(\pk_s8ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[10]  ( .Q(\pk_s9ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[5]  ( .Q(\pk_saba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[15]  ( .Q(\pk_sbba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[4]  ( .Q(\pk_scba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[15]  ( .Q(\pk_sfba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[7]  ( .Q(\pk_saba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[17]  ( .Q(\pk_sbba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[13]  ( .Q(\pk_sdba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[2]  ( .Q(\pk_s3ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[12]  ( .Q(\pk_s9ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[11]  ( .Q(\pk_sdba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[8]  ( .Q(\pk_sdba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[9]  ( .Q(\pk_sfba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[6]  ( .Q(\pk_scba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[17]  ( .Q(\pk_sfba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff51/U839  ( .ZN(\REGF/pbmemff51/n4469 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_invx2 \REGF/pbmemff51/U844  ( .ZN(\REGF/pbmemff51/n4477 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[16]  ( .Q(\pk_s0ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[12]  ( .Q(\pk_s0ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[14]  ( .Q(\pk_s2ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[12]  ( .Q(\pk_s4ba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[3]  ( .Q(\pk_s8ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[0]  ( .Q(\pk_sfba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[5]  ( .Q(\pk_s4ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[14]  ( .Q(\pk_s6ba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[4]  ( .Q(\pk_s6ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[7]  ( .Q(\pk_s1ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[6]  ( .Q(\pk_s3ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[9]  ( .Q(\pk_s6ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[18]  ( .Q(
        \REGF/pk_sdba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[1]  ( .Q(\pk_sdba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[13]  ( .Q(\pk_sfba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[2]  ( .Q(\pk_scba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[16]  ( .Q(\pk_s9ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[15]  ( .Q(\pk_sdba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[8]  ( .Q(\pk_s4ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[3]  ( .Q(\pk_saba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[13]  ( .Q(\pk_sbba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[10]  ( .Q(\pk_s2ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[1]  ( .Q(\pk_s4ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[10]  ( .Q(\pk_s6ba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SDBA19B_reg[5]  ( .Q(\pk_sdba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[22] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S6BA19B_reg[0]  ( .Q(\pk_s6ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[29] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S4BA19B_reg[16]  ( .Q(\pk_s4ba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[31] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SFBA19B_reg[4]  ( .Q(\pk_sfba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[20] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[3]  ( .Q(\pk_s2ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[18]  ( .Q(
        \REGF/pk_s3ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[4]  ( .Q(\pk_s5ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[7]  ( .Q(\pk_s8ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[14]  ( .Q(\pk_seba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[0]  ( .Q(\pk_seba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[18]  ( .Q(
        \REGF/pk_s7ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[12]  ( .Q(\pk_scba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[11]  ( .Q(\pk_s3ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[5]  ( .Q(\pk_s7ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[17]  ( .Q(\pk_s8ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[2]  ( .Q(\pk_s9ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[14]  ( .Q(\pk_saba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[7]  ( .Q(\pk_sbba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[17]  ( .Q(\pk_s5ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_invx1 \REGF/pbmemff51/U845  ( .ZN(\REGF/pbmemff51/n4473 ), .A(
        \REGF/n8052 ) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[2]  ( .Q(\pk_s0ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[9]  ( .Q(\pk_seba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[17]  ( .Q(\pk_s1ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[11]  ( .Q(\pk_s7ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[1]  ( .Q(\pk_s7ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[13]  ( .Q(\pk_s8ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[6]  ( .Q(\pk_s9ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[10]  ( .Q(\pk_saba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[6]  ( .Q(\pk_s0ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[9]  ( .Q(\pk_s5ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[0]  ( .Q(\pk_s5ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[16]  ( .Q(\pk_scba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[10]  ( .Q(\pk_seba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[4]  ( .Q(\pk_seba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[15]  ( .Q(\pk_s7ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[4]  ( .Q(\pk_s0ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[13]  ( .Q(\pk_s1ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[7]  ( .Q(\pk_s2ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[13]  ( .Q(\pk_s5ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[5]  ( .Q(\pk_s2ba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[15]  ( .Q(\pk_s3ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[3]  ( .Q(\pk_sbba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[8]  ( .Q(\pk_s7ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[18]  ( .Q(
        \REGF/pk_s8ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[17]  ( .Q(\pk_s3ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[11]  ( .Q(\pk_s5ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[17]  ( .Q(\pk_s7ba_h[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4471 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[1]  ( .Q(\pk_sbba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[11]  ( .Q(\pk_s1ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_invx2 \REGF/pbmemff51/U842  ( .ZN(\REGF/pbmemff51/n4471 ), .A(
        \REGF/pbmemff51/n4473 ) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[18]  ( .Q(
        \REGF/pk_s1ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[2]  ( .Q(\pk_s5ba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[14]  ( .Q(\pk_scba_h[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[6]  ( .Q(\pk_seba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[18]  ( .Q(
        \REGF/pk_s5ba_h[18] ), .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 
        ), .SD(PDLIN[18]), .SE(\pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[4]  ( .Q(\pk_s9ba_h[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[12]  ( .Q(\pk_seba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[3]  ( .Q(\pk_s7ba_h[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[11]  ( .Q(\pk_s8ba_h[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4475 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[12]  ( .Q(\pk_saba_h[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[9]  ( .Q(\pk_s0ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S0BA19B_reg[0]  ( .Q(\pk_s0ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[35] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[8]  ( .Q(\pk_sbba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S1BA19B_reg[15]  ( .Q(\pk_s1ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[34] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[8]  ( .Q(\pk_s2ba_h[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S2BA19B_reg[1]  ( .Q(\pk_s2ba_h[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[33] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S3BA19B_reg[13]  ( .Q(\pk_s3ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[32] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[13]  ( .Q(\pk_s7ba_h[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SBBA19B_reg[5]  ( .Q(\pk_sbba_h[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[24] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[15]  ( .Q(\pk_s5ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S7BA19B_reg[7]  ( .Q(\pk_s7ba_h[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[28] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[9]  ( .Q(\pk_s9ba_h[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S8BA19B_reg[15]  ( .Q(\pk_s8ba_h[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4476 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[27] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S9BA19B_reg[0]  ( .Q(\pk_s9ba_h[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4474 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[26] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SABA19B_reg[16]  ( .Q(\pk_saba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[25] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[16]  ( .Q(\pk_seba_h[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4472 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_S5BA19B_reg[6]  ( .Q(\pk_s5ba_h[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4469 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[30] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SEBA19B_reg[2]  ( .Q(\pk_seba_h[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4470 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[21] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff51/RO_SCBA19B_reg[10]  ( .Q(\pk_scba_h[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff51/n4477 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[23] ), .CP(SCLK) );
    snl_ao222x1 \UPIF/CSGN/U1468  ( .Z(\pk_rwrit_h[52] ), .A(\pk_rread_h[44] ), 
        .B(\UPIF/reg_wr ), .C(ph_srcadr1_h), .D(\UPIF/CSGN/n1694 ), .E(
        ph_oprtrs_h), .F(st_exectl) );
    snl_and23x1 \UPIF/CSGN/U1474  ( .Z(\UPIF/CSGN/n1724 ), .A(
        \UPIF/CSGN/n1725 ), .B(PA[3]), .C(PA[5]) );
    snl_nor02x2 \UPIF/CSGN/U1483  ( .ZN(\pk_rwrit_h[12] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1708 ) );
    snl_and02x2 \UPIF/CSGN/U1498  ( .Z(\pk_rread_h[43] ), .A(\UPIF/CSGN/n1747 
        ), .B(\UPIF/CSGN/n1736 ) );
    snl_nor02x3 \UPIF/CSGN/U1508  ( .ZN(\pk_rwrit_h[39] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1660 ) );
    snl_invx2 \UPIF/CSGN/U1541  ( .ZN(\pk_rread_h[4] ), .A(\UPIF/CSGN/n1709 )
         );
    snl_invx2 \UPIF/CSGN/U1566  ( .ZN(\pk_rread_h[30] ), .A(\UPIF/CSGN/n1686 )
         );
    snl_nand02x1 \UPIF/CSGN/U1656  ( .ZN(\UPIF/CSGN/n1662 ), .A(
        \UPIF/CSGN/n1742 ), .B(\UPIF/CSGN/n1736 ) );
    snl_nand03x0 \UPIF/CSGN/U1638  ( .ZN(\UPIF/CSGN/n1654 ), .A(
        \UPIF/CSGN/n1729 ), .B(PA[6]), .C(PA[7]) );
    snl_nand02x1 \UPIF/CSGN/U1671  ( .ZN(\UPIF/CSGN/n1695 ), .A(
        \UPIF/CSGN/n1747 ), .B(\UPIF/CSGN/n1740 ) );
    snl_nor02x3 \UPIF/CSGN/U1513  ( .ZN(\pk_rwrit_h[40] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1668 ) );
    snl_and02x1 \UPIF/CSGN/U1583  ( .Z(\pk_rwrit_h[21] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[14] ) );
    snl_nand02x1 \UPIF/CSGN/U1694  ( .ZN(\UPIF/CSGN/n1681 ), .A(
        \UPIF/CSGN/n1756 ), .B(\UPIF/CSGN/n1728 ) );
    snl_nand12x1 \UPIF/CSGN/U1704  ( .ZN(\UPIF/CSGN/n1758 ), .A(
        \UPIF/CSGN/n1718 ), .B(PA[11]) );
    snl_invx05 \UPIF/CSGN/U1723  ( .ZN(\UPIF/CSGN/n1728 ), .A(
        \UPIF/CSGN/n1676 ) );
    snl_oai013x0 \UPIF/CSGN/U1598  ( .ZN(cnt_write_h), .A(\UPIF/CSGN/n1639 ), 
        .B(\UPIF/CSGN/n1679 ), .C(\UPIF/CSGN/n1676 ), .D(\UPIF/CSGN/n1680 ) );
    snl_invx05 \UPIF/CSGN/U1738  ( .ZN(\UPIF/CSGN/reg_stat_h ), .A(
        \UPIF/CSGN/n1758 ) );
    snl_invx2 \UPIF/CSGN/U1534  ( .ZN(\pk_rread_h[52] ), .A(\UPIF/CSGN/n1703 )
         );
    snl_and02x1 \UPIF/CSGN/U1604  ( .Z(\pk_rwrit_h[11] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[11] ) );
    snl_nand02x1 \UPIF/CSGN/U1623  ( .ZN(\UPIF/CSGN/n1679 ), .A(PA[6]), .B(
        \UPIF/CSGN/n1723 ) );
    snl_nor02x2 \UPIF/CSGN/U1491  ( .ZN(\pk_rwrit_h[28] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1656 ) );
    snl_invx2 \UPIF/CSGN/U1548  ( .ZN(\pk_rread_h[27] ), .A(\UPIF/CSGN/n1667 )
         );
    snl_nand02x1 \UPIF/CSGN/U1678  ( .ZN(\UPIF/CSGN/n1677 ), .A(
        \UPIF/CSGN/n1733 ), .B(\UPIF/CSGN/n1732 ) );
    snl_and02x2 \UPIF/CSGN/U1501  ( .Z(\pk_rread_h[42] ), .A(\UPIF/CSGN/n1748 
        ), .B(\UPIF/CSGN/n1736 ) );
    snl_nor02x3 \UPIF/CSGN/U1526  ( .ZN(\pk_rread_h[46] ), .A(
        \UPIF/CSGN/n1683 ), .B(\UPIF/CSGN/n1689 ) );
    snl_nor02x1 \UPIF/CSGN/U1616  ( .ZN(\pk_rwrit_h[4] ), .A(\UPIF/CSGN/n1639 
        ), .B(\UPIF/CSGN/n1709 ) );
    snl_nand03x0 \UPIF/CSGN/U1631  ( .ZN(\UPIF/CSGN/n1665 ), .A(
        \UPIF/CSGN/n1729 ), .B(\UPIF/CSGN/n1649 ), .C(PA[7]) );
    snl_invx2 \UPIF/CSGN/U1553  ( .ZN(\pk_rread_h[49] ), .A(\UPIF/CSGN/n1641 )
         );
    snl_nand04x0 \UPIF/CSGN/U1574  ( .ZN(\UPIF/CSGN/*cell*4224/U3/CONTROL1 ), 
        .A(\UPIF/CSGN/n1640 ), .B(\UPIF/CSGN/n1641 ), .C(\UPIF/CSGN/n1642 ), 
        .D(\UPIF/CSGN/n1643 ) );
    snl_nor03x0 \UPIF/CSGN/U1591  ( .ZN(\UPIF/CSGN/n_1054 ), .A(
        \UPIF/CSGN/n1643 ), .B(WR), .C(\UPIF/CSGN/n1642 ) );
    snl_nand02x1 \UPIF/CSGN/U1686  ( .ZN(\UPIF/CSGN/n1678 ), .A(
        \UPIF/CSGN/n1750 ), .B(\UPIF/CSGN/n1724 ) );
    snl_aoi022x1 \UPIF/CSGN/U1716  ( .ZN(\UPIF/CSGN/n1712 ), .A(po_imdselh), 
        .B(st_exectl), .C(\pk_rread_h[42] ), .D(\UPIF/reg_wr ) );
    snl_invx05 \UPIF/CSGN/U1731  ( .ZN(\UPIF/CSGN/n1670 ), .A(
        \UPIF/CSGN/n1757 ) );
    snl_nand02x1 \UPIF/CSGN/U1644  ( .ZN(\UPIF/CSGN/n1690 ), .A(
        \UPIF/CSGN/n1734 ), .B(\UPIF/CSGN/n1731 ) );
    snl_invx2 \UPIF/CSGN/U1554  ( .ZN(\pk_rread_h[21] ), .A(\UPIF/CSGN/n1656 )
         );
    snl_nand02x1 \UPIF/CSGN/U1663  ( .ZN(\UPIF/CSGN/n1703 ), .A(
        \UPIF/CSGN/n1744 ), .B(\UPIF/CSGN/n1738 ) );
    snl_nand02x1 \UPIF/CSGN/U1664  ( .ZN(\UPIF/CSGN/n1692 ), .A(
        \UPIF/CSGN/n1743 ), .B(\UPIF/CSGN/n1741 ) );
    snl_invx2 \UPIF/CSGN/U1573  ( .ZN(\pk_rread_h[38] ), .A(\UPIF/CSGN/n1702 )
         );
    snl_nand02x1 \UPIF/CSGN/U1643  ( .ZN(\UPIF/CSGN/n1698 ), .A(
        \UPIF/CSGN/n1733 ), .B(\UPIF/CSGN/n1728 ) );
    snl_ao222x2 \UPIF/CSGN/U1469  ( .Z(\pk_rwrit_h[66] ), .A(\pk_rread_h[61] ), 
        .B(\UPIF/reg_wr ), .C(ph_dprtrs_h), .D(\UPIF/CSGN/n1694 ), .E(
        st_exectl), .F(wdpr) );
    snl_invx1 \UPIF/CSGN/U1472  ( .ZN(\UPIF/CSGN/n1639 ), .A(\UPIF/reg_wr ) );
    snl_invx2 \UPIF/CSGN/U1473  ( .ZN(\UPIF/CSGN/n1650 ), .A(\UPIF/reg_wr ) );
    snl_nor02x2 \UPIF/CSGN/U1496  ( .ZN(\pk_rwrit_h[24] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1693 ) );
    snl_nor02x3 \UPIF/CSGN/U1506  ( .ZN(\pk_rwrit_h[36] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1657 ) );
    snl_nor02x3 \UPIF/CSGN/U1521  ( .ZN(\pk_rread_h[37] ), .A(
        \UPIF/CSGN/n1688 ), .B(\UPIF/CSGN/n1646 ) );
    snl_and02x1 \UPIF/CSGN/U1596  ( .Z(\pk_rwrit_h[20] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[13] ) );
    snl_nand02x1 \UPIF/CSGN/U1681  ( .ZN(\UPIF/CSGN/n1660 ), .A(
        \UPIF/CSGN/n1750 ), .B(\UPIF/CSGN/n1734 ) );
    snl_nor04x0 \UPIF/CSGN/U1711  ( .ZN(\UPIF/CSGN/n1717 ), .A(PA[22]), .B(PA
        [23]), .C(PA[24]), .D(PA[25]) );
    snl_or02x1 \UPIF/CSGN/U1736  ( .Z(\UPIF/CSGN/n1715 ), .A(ph_sprlth), .B(
        \UPIF/CSGN/n1638 ) );
    snl_nor02x1 \UPIF/CSGN/U1611  ( .ZN(\pk_rwrit_h[48] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1701 ) );
    snl_nand12x1 \UPIF/CSGN/U1636  ( .ZN(\UPIF/CSGN/n1652 ), .A(
        \UPIF/CSGN/n1679 ), .B(\UPIF/CSGN/n1724 ) );
    snl_nor02x2 \UPIF/CSGN/U1484  ( .ZN(\pk_rwrit_h[32] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1691 ) );
    snl_invx2 \UPIF/CSGN/U1533  ( .ZN(\pk_rread_h[48] ), .A(\UPIF/CSGN/n1685 )
         );
    snl_invx2 \UPIF/CSGN/U1568  ( .ZN(\pk_rread_h[58] ), .A(\UPIF/CSGN/n1662 )
         );
    snl_nand02x1 \UPIF/CSGN/U1658  ( .ZN(\UPIF/CSGN/n1651 ), .A(
        \UPIF/CSGN/n1742 ), .B(\UPIF/CSGN/n1740 ) );
    snl_nand02x1 \UPIF/CSGN/U1688  ( .ZN(\UPIF/CSGN/n1696 ), .A(PA[4]), .B(
        \UPIF/CSGN/n1724 ) );
    snl_invx05 \UPIF/CSGN/U1718  ( .ZN(ret_cont_h), .A(\UPIF/CSGN/n1659 ) );
    snl_nor03x0 \UPIF/CSGN/U1603  ( .ZN(ph_schvx_h), .A(\UPIF/CSGN/n1688 ), 
        .B(\UPIF/CSGN/n1639 ), .C(\UPIF/CSGN/n1689 ) );
    snl_nor02x1 \UPIF/CSGN/U1624  ( .ZN(\UPIF/CSGN/n1726 ), .A(
        \UPIF/CSGN/n1725 ), .B(PA[5]) );
    snl_nor02x3 \UPIF/CSGN/U1514  ( .ZN(\pk_rwrit_h[43] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1706 ) );
    snl_invx1 \UPIF/CSGN/U1528  ( .ZN(\pk_rwrit_h[59] ), .A(\UPIF/CSGN/n1680 )
         );
    snl_or08x1 \UPIF/CSGN/U1618  ( .Z(\UPIF/CSGN/n1718 ), .A(PA[15]), .B(PA
        [16]), .C(PA[12]), .D(PA[14]), .E(PA[17]), .F(PA[18]), .G(PA[19]), .H(
        \UPIF/CSGN/n1719 ) );
    snl_invx2 \UPIF/CSGN/U1546  ( .ZN(\pk_rread_h[3] ), .A(\UPIF/CSGN/n1677 )
         );
    snl_nor02x1 \UPIF/CSGN/U1584  ( .ZN(\pk_rwrit_h[60] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1663 ) );
    snl_nand02x1 \UPIF/CSGN/U1676  ( .ZN(\UPIF/CSGN/n1655 ), .A(
        \UPIF/CSGN/n1747 ), .B(\UPIF/CSGN/n1744 ) );
    snl_nand02x1 \UPIF/CSGN/U1693  ( .ZN(\UPIF/CSGN/n1697 ), .A(
        \UPIF/CSGN/n1756 ), .B(\UPIF/CSGN/n1734 ) );
    snl_invx05 \UPIF/CSGN/U1724  ( .ZN(\UPIF/CSGN/n1734 ), .A(
        \UPIF/CSGN/n1671 ) );
    snl_nand02x1 \UPIF/CSGN/U1703  ( .ZN(\UPIF/CSGN/n1708 ), .A(
        \UPIF/CSGN/n1757 ), .B(\UPIF/CSGN/n1724 ) );
    snl_invx2 \UPIF/CSGN/U1561  ( .ZN(\pk_rread_h[17] ), .A(\UPIF/CSGN/n1693 )
         );
    snl_and02x1 \UPIF/CSGN/U1651  ( .Z(\UPIF/CSGN/n1739 ), .A(
        \UPIF/CSGN/n1735 ), .B(PA[4]) );
    snl_and02x2 \UPIF/CSGN/U1497  ( .Z(\pk_rread_h[45] ), .A(\UPIF/CSGN/n1745 
        ), .B(\UPIF/CSGN/n1740 ) );
    snl_nor02x3 \UPIF/CSGN/U1520  ( .ZN(\pk_rread_h[1] ), .A(\UPIF/CSGN/n1671 
        ), .B(\UPIF/CSGN/n1679 ) );
    snl_invx2 \UPIF/CSGN/U1569  ( .ZN(\pk_rread_h[18] ), .A(\UPIF/CSGN/n1682 )
         );
    snl_and23x0 \UPIF/CSGN/U1659  ( .Z(\UPIF/CSGN/n1743 ), .A(
        \UPIF/CSGN/n1649 ), .B(PA[4]), .C(\UPIF/CSGN/n1735 ) );
    snl_nor03x0 \UPIF/CSGN/U1610  ( .ZN(\pk_rwrit_h[19] ), .A(
        \UPIF/CSGN/n1699 ), .B(\UPIF/CSGN/n1700 ), .C(\UPIF/CSGN/n1639 ) );
    snl_nand03x0 \UPIF/CSGN/U1637  ( .ZN(\UPIF/CSGN/n1699 ), .A(PA[5]), .B(
        \UPIF/CSGN/n1720 ), .C(PA[3]) );
    snl_nor02x3 \UPIF/CSGN/U1507  ( .ZN(\pk_rwrit_h[38] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1710 ) );
    snl_invx2 \UPIF/CSGN/U1555  ( .ZN(\pk_rread_h[57] ), .A(\UPIF/CSGN/n1675 )
         );
    snl_nor03x0 \UPIF/CSGN/U1597  ( .ZN(\pk_rwrit_h[13] ), .A(
        \UPIF/CSGN/n1654 ), .B(\UPIF/CSGN/n1647 ), .C(\UPIF/CSGN/n1639 ) );
    snl_nand02x1 \UPIF/CSGN/U1665  ( .ZN(\UPIF/CSGN/n1683 ), .A(PA[7]), .B(
        \UPIF/CSGN/n1728 ) );
    snl_and02x1 \UPIF/CSGN/U1680  ( .Z(\UPIF/CSGN/n1750 ), .A(
        \UPIF/CSGN/n1749 ), .B(\UPIF/CSGN/n1727 ) );
    snl_invx05 \UPIF/CSGN/U1737  ( .ZN(\UPIF/CSGN/n1725 ), .A(
        \UPIF/CSGN/n1720 ) );
    snl_nor02x1 \UPIF/CSGN/U1710  ( .ZN(\UPIF/CSGN/n1640 ), .A(
        \pk_rread_h[50] ), .B(\pk_rread_h[47] ) );
    snl_invx2 \UPIF/CSGN/U1572  ( .ZN(\pk_rread_h[63] ), .A(\UPIF/CSGN/n1714 )
         );
    snl_nand02x1 \UPIF/CSGN/U1642  ( .ZN(\UPIF/CSGN/n1669 ), .A(
        \UPIF/CSGN/n1734 ), .B(\UPIF/CSGN/n1733 ) );
    snl_ao223x2 \UPIF/CSGN/U1470  ( .Z(\pk_rwrit_h[65] ), .A(ph_adrwtenh), .B(
        \UPIF/CSGN/n1715 ), .C(ph_sprtrs_h), .D(\pk_rread_h[60] ), .E(
        \UPIF/reg_wr ), .F(wspr), .G(st_exectl) );
    snl_and34x1 \UPIF/CSGN/U1475  ( .Z(code_area_h), .A(PA[27]), .B(PA[29]), 
        .C(\UPIF/CSGN/n1644 ), .D(PA[28]) );
    snl_nor02x2 \UPIF/CSGN/U1482  ( .ZN(\pk_rwrit_h[26] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1705 ) );
    snl_and02x2 \UPIF/CSGN/U1485  ( .Z(\pk_rread_h[44] ), .A(\UPIF/CSGN/n1746 
        ), .B(\UPIF/CSGN/n1740 ) );
    snl_nor02x3 \UPIF/CSGN/U1515  ( .ZN(\pk_rwrit_h[42] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1673 ) );
    snl_oai023x2 \UPIF/CSGN/U1529  ( .ZN(\pk_rwrit_h[68] ), .A(
        \UPIF/CSGN/n1713 ), .B(phsaerrh), .C(\UPIF/alusfterr ), .D(
        \UPIF/CSGN/n1639 ), .E(\UPIF/CSGN/n1714 ) );
    snl_invx2 \UPIF/CSGN/U1547  ( .ZN(\pk_rread_h[7] ), .A(\UPIF/CSGN/n1698 )
         );
    snl_nand02x1 \UPIF/CSGN/U1677  ( .ZN(\UPIF/CSGN/n1668 ), .A(
        \UPIF/CSGN/n1748 ), .B(\UPIF/CSGN/n1744 ) );
    snl_invx2 \UPIF/CSGN/U1560  ( .ZN(\pk_rread_h[5] ), .A(\UPIF/CSGN/n1687 )
         );
    snl_nor02x1 \UPIF/CSGN/U1619  ( .ZN(\UPIF/CSGN/n1720 ), .A(
        \UPIF/CSGN/n1718 ), .B(PA[11]) );
    snl_and02x1 \UPIF/CSGN/U1650  ( .Z(\UPIF/CSGN/n1694 ), .A(
        \UPIF/CSGN/n1638 ), .B(ph_adrwtenh) );
    snl_invx2 \UPIF/CSGN/U1532  ( .ZN(\pk_rread_h[56] ), .A(\UPIF/CSGN/n1651 )
         );
    snl_nor03x0 \UPIF/CSGN/U1585  ( .ZN(\pk_rwrit_h[17] ), .A(
        \UPIF/CSGN/n1664 ), .B(\UPIF/CSGN/n1665 ), .C(\UPIF/CSGN/n1639 ) );
    snl_nand02x1 \UPIF/CSGN/U1689  ( .ZN(\UPIF/CSGN/n1661 ), .A(
        \UPIF/CSGN/n1753 ), .B(\UPIF/CSGN/n1749 ) );
    snl_and02x1 \UPIF/CSGN/U1692  ( .Z(\UPIF/CSGN/n1756 ), .A(
        \UPIF/CSGN/n1755 ), .B(\UPIF/CSGN/n1727 ) );
    snl_nor02x1 \UPIF/CSGN/U1702  ( .ZN(\UPIF/CSGN/n1757 ), .A(
        \UPIF/CSGN/n1654 ), .B(PA[4]) );
    snl_invx05 \UPIF/CSGN/U1725  ( .ZN(\UPIF/CSGN/n1736 ), .A(
        \UPIF/CSGN/n1689 ) );
    snl_invx05 \UPIF/CSGN/U1719  ( .ZN(write_pr_h), .A(\UPIF/CSGN/n1652 ) );
    snl_nor02x1 \UPIF/CSGN/U1602  ( .ZN(\pk_rwrit_h[5] ), .A(\UPIF/CSGN/n1650 
        ), .B(\UPIF/CSGN/n1687 ) );
    snl_nand02x1 \UPIF/CSGN/U1625  ( .ZN(\UPIF/CSGN/n1676 ), .A(PA[3]), .B(
        \UPIF/CSGN/n1726 ) );
    snl_nor03x0 \UPIF/CSGN/U1599  ( .ZN(\pk_rwrit_h[44] ), .A(
        \UPIF/CSGN/n1683 ), .B(\UPIF/CSGN/n1639 ), .C(\UPIF/CSGN/n1646 ) );
    snl_sffqrnx1 \UPIF/CSGN/err_fact_w_reg  ( .Q(\pk_rwrit_h[0] ), .D(1'b0), 
        .RN(n10733), .SD(\UPIF/CSGN/*cell*4224/U3/CONTROL1 ), .SE(
        \UPIF/CSGN/n_1054 ), .CP(SCLK) );
    snl_nor02x2 \UPIF/CSGN/U1490  ( .ZN(\pk_rwrit_h[30] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1681 ) );
    snl_and02x2 \UPIF/CSGN/U1499  ( .Z(\pk_rread_h[61] ), .A(\UPIF/CSGN/n1740 
        ), .B(\UPIF/CSGN/n1737 ) );
    snl_nor02x3 \UPIF/CSGN/U1512  ( .ZN(\pk_rwrit_h[58] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1703 ) );
    snl_invx2 \UPIF/CSGN/U1535  ( .ZN(\pk_rread_h[20] ), .A(\UPIF/CSGN/n1674 )
         );
    snl_nor02x1 \UPIF/CSGN/U1605  ( .ZN(\pk_rwrit_h[57] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1692 ) );
    snl_invx05 \UPIF/CSGN/U1622  ( .ZN(\UPIF/CSGN/n1649 ), .A(PA[6]) );
    snl_nand02x1 \UPIF/CSGN/U1639  ( .ZN(\UPIF/CSGN/n1664 ), .A(
        \UPIF/CSGN/n1732 ), .B(PA[4]) );
    snl_and02x2 \UPIF/CSGN/U1500  ( .Z(\pk_rread_h[62] ), .A(\UPIF/CSGN/n1738 
        ), .B(\UPIF/CSGN/n1736 ) );
    snl_nor02x3 \UPIF/CSGN/U1509  ( .ZN(\pk_rwrit_h[7] ), .A(\UPIF/CSGN/n1650 
        ), .B(\UPIF/CSGN/n1698 ) );
    snl_invx2 \UPIF/CSGN/U1540  ( .ZN(\pk_rread_h[28] ), .A(\UPIF/CSGN/n1678 )
         );
    snl_invx2 \UPIF/CSGN/U1567  ( .ZN(\pk_rread_h[22] ), .A(\UPIF/CSGN/n1707 )
         );
    snl_and02x1 \UPIF/CSGN/U1582  ( .Z(\pk_rwrit_h[1] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[1] ) );
    snl_nand02x1 \UPIF/CSGN/U1695  ( .ZN(\UPIF/CSGN/n1672 ), .A(
        \UPIF/CSGN/n1732 ), .B(\UPIF/CSGN/n1731 ) );
    snl_invx05 \UPIF/CSGN/U1705  ( .ZN(\UPIF/CSGN/n1684 ), .A(
        \UPIF/tr_count_lt ) );
    snl_invx05 \UPIF/CSGN/U1722  ( .ZN(\UPIF/CSGN/n1732 ), .A(
        \UPIF/CSGN/n1699 ) );
    snl_nand02x1 \UPIF/CSGN/U1657  ( .ZN(\UPIF/CSGN/n1675 ), .A(
        \UPIF/CSGN/n1741 ), .B(\UPIF/CSGN/n1740 ) );
    snl_sffqrnx1 \UPIF/CSGN/pk_rwrit56h_reg  ( .Q(\pk_rwrit_h[56] ), .D(1'b0), 
        .RN(n10733), .SD(\UPIF/CSGN/*cell*4224/U3/CONTROL1 ), .SE(
        \UPIF/CSGN/n_1040 ), .CP(SCLK) );
    snl_invx2 \UPIF/CSGN/U1552  ( .ZN(\pk_rread_h[23] ), .A(\UPIF/CSGN/n1681 )
         );
    snl_nor03x0 \UPIF/CSGN/U1575  ( .ZN(\UPIF/write_by_h ), .A(
        \UPIF/CSGN/n1647 ), .B(\UPIF/CSGN/n1648 ), .C(\UPIF/CSGN/n1649 ) );
    snl_nor03x0 \UPIF/CSGN/U1645  ( .ZN(\UPIF/CSGN/n1735 ), .A(PA[8]), .B(PA
        [10]), .C(PA[9]) );
    snl_nand02x1 \UPIF/CSGN/U1670  ( .ZN(\UPIF/CSGN/n1709 ), .A(
        \UPIF/CSGN/n1733 ), .B(\UPIF/CSGN/n1724 ) );
    snl_ao012x1 \UPIF/CSGN/U1590  ( .Z(\pk_rwrit_h[54] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[46] ), .C(ph_stregwt_h) );
    snl_nand02x1 \UPIF/CSGN/U1662  ( .ZN(\UPIF/CSGN/n1646 ), .A(
        \UPIF/CSGN/n1739 ), .B(PA[6]) );
    snl_nand02x1 \UPIF/CSGN/U1687  ( .ZN(\UPIF/CSGN/n1667 ), .A(
        \UPIF/CSGN/n1750 ), .B(\UPIF/CSGN/n1732 ) );
    snl_invx05 \UPIF/CSGN/U1717  ( .ZN(\UPIF/CSGN/n1643 ), .A(\pk_rread_h[0] )
         );
    snl_invx05 \UPIF/CSGN/U1730  ( .ZN(\UPIF/CSGN/n1754 ), .A(
        \UPIF/CSGN/n1664 ) );
    snl_nor02x3 \UPIF/CSGN/U1527  ( .ZN(\pk_rread_h[50] ), .A(PA[10]), .B(
        \UPIF/CSGN/n1758 ) );
    snl_nand02x1 \UPIF/CSGN/U1617  ( .ZN(\UPIF/CSGN/n1644 ), .A(
        \UPIF/CSGN/n1716 ), .B(\UPIF/CSGN/n1717 ) );
    snl_invx05 \UPIF/CSGN/U1630  ( .ZN(\UPIF/CSGN/n1722 ), .A(PA[7]) );
    snl_and02x2 \UPIF/CSGN/U1477  ( .Z(\pk_rwrit_h[9] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[9] ) );
    snl_nor02x2 \UPIF/CSGN/U1480  ( .ZN(\pk_rwrit_h[27] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1674 ) );
    snl_invx2 \UPIF/CSGN/U1537  ( .ZN(\pk_rread_h[24] ), .A(\UPIF/CSGN/n1697 )
         );
    snl_invx2 \UPIF/CSGN/U1542  ( .ZN(\pk_rread_h[8] ), .A(\UPIF/CSGN/n1669 )
         );
    snl_invx2 \UPIF/CSGN/U1549  ( .ZN(\pk_rread_h[59] ), .A(\UPIF/CSGN/n1666 )
         );
    snl_and23x0 \UPIF/CSGN/U1679  ( .Z(\UPIF/CSGN/n1749 ), .A(PA[7]), .B(PA[6]
        ), .C(\UPIF/CSGN/n1729 ) );
    snl_invx2 \UPIF/CSGN/U1565  ( .ZN(\pk_rread_h[26] ), .A(\UPIF/CSGN/n1661 )
         );
    snl_nor02x1 \UPIF/CSGN/U1655  ( .ZN(\UPIF/CSGN/n1742 ), .A(
        \UPIF/CSGN/n1699 ), .B(PA[7]) );
    snl_nand02x1 \UPIF/CSGN/U1672  ( .ZN(\UPIF/CSGN/n1701 ), .A(
        \UPIF/CSGN/n1748 ), .B(\UPIF/CSGN/n1740 ) );
    snl_nor02x1 \UPIF/CSGN/U1580  ( .ZN(\UPIF/CSGN/n_1040 ), .A(
        \UPIF/CSGN/n1640 ), .B(\UPIF/CSGN/n1642 ) );
    snl_invx05 \UPIF/CSGN/U1720  ( .ZN(\UPIF/CSGN/n1704 ), .A(\UPIF/alusfterr 
        ) );
    snl_ao022x1 \UPIF/CSGN/U1607  ( .Z(\pk_rwrit_h[51] ), .A(\pk_rread_h[43] ), 
        .B(\UPIF/reg_wr ), .C(ph_srcadr2_h), .D(\UPIF/CSGN/n1694 ) );
    snl_nand02x1 \UPIF/CSGN/U1697  ( .ZN(\UPIF/CSGN/n1656 ), .A(
        \UPIF/CSGN/n1755 ), .B(\UPIF/CSGN/n1752 ) );
    snl_invx05 \UPIF/CSGN/U1707  ( .ZN(\UPIF/CSGN/n1642 ), .A(\UPIF/ready_eoc 
        ) );
    snl_nor02x3 \UPIF/CSGN/U1510  ( .ZN(\pk_rwrit_h[41] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1655 ) );
    snl_invx2 \UPIF/CSGN/U1559  ( .ZN(\pk_rread_h[29] ), .A(\UPIF/CSGN/n1657 )
         );
    snl_nand14x0 \UPIF/CSGN/U1620  ( .ZN(\UPIF/CSGN/n1648 ), .A(PA[10]), .B(PA
        [9]), .C(\UPIF/CSGN/n1721 ), .D(\UPIF/CSGN/n1722 ) );
    snl_nor02x1 \UPIF/CSGN/U1669  ( .ZN(\UPIF/CSGN/n1748 ), .A(
        \UPIF/CSGN/n1699 ), .B(\UPIF/CSGN/n1722 ) );
    snl_sffqrnx1 \UPIF/CSGN/ex_stat1_w_reg  ( .Q(\pk_rwrit_h[55] ), .D(1'b0), 
        .RN(n10733), .SD(\UPIF/CSGN/*cell*4224/U3/CONTROL1 ), .SE(
        \UPIF/CSGN/n_1047 ), .CP(SCLK) );
    snl_nor02x2 \UPIF/CSGN/U1489  ( .ZN(\pk_rwrit_h[31] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1697 ) );
    snl_nor02x2 \UPIF/CSGN/U1492  ( .ZN(\pk_rwrit_h[29] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1707 ) );
    snl_nor02x2 \UPIF/CSGN/U1502  ( .ZN(\pk_rwrit_h[2] ), .A(\UPIF/CSGN/n1650 
        ), .B(\UPIF/CSGN/n1672 ) );
    snl_nor02x3 \UPIF/CSGN/U1525  ( .ZN(\pk_rread_h[13] ), .A(
        \UPIF/CSGN/n1665 ), .B(\UPIF/CSGN/n1647 ) );
    snl_ao012x1 \UPIF/CSGN/U1589  ( .Z(\pk_rwrit_h[47] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[39] ), .C(phsaerrh) );
    snl_nor02x1 \UPIF/CSGN/U1615  ( .ZN(ph_sastlth), .A(\UPIF/CSGN/n1701 ), 
        .B(\UPIF/CSGN/n1684 ) );
    snl_invx05 \UPIF/CSGN/U1729  ( .ZN(\UPIF/CSGN/n1753 ), .A(
        \UPIF/CSGN/n1696 ) );
    snl_nor02x3 \UPIF/CSGN/U1519  ( .ZN(\pk_rread_h[11] ), .A(
        \UPIF/CSGN/n1670 ), .B(\UPIF/CSGN/n1699 ) );
    snl_nor03x0 \UPIF/CSGN/U1629  ( .ZN(\UPIF/CSGN/n1729 ), .A(PA[9]), .B(PA
        [10]), .C(\UPIF/CSGN/n1721 ) );
    snl_nor02x1 \UPIF/CSGN/U1632  ( .ZN(\UPIF/CSGN/n1730 ), .A(
        \UPIF/CSGN/n1665 ), .B(PA[4]) );
    snl_nor02x2 \UPIF/CSGN/U1495  ( .ZN(\pk_rwrit_h[35] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1678 ) );
    snl_invx2 \UPIF/CSGN/U1539  ( .ZN(\pk_rread_h[36] ), .A(\UPIF/CSGN/n1706 )
         );
    snl_invx2 \UPIF/CSGN/U1550  ( .ZN(\pk_rread_h[19] ), .A(\UPIF/CSGN/n1705 )
         );
    snl_nor02x1 \UPIF/CSGN/U1592  ( .ZN(\pk_rwrit_h[62] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1675 ) );
    snl_invx05 \UPIF/CSGN/U1732  ( .ZN(\UPIF/CSGN/n1700 ), .A(
        \UPIF/CSGN/n1730 ) );
    snl_nand02x1 \UPIF/CSGN/U1685  ( .ZN(\UPIF/CSGN/n1657 ), .A(
        \UPIF/CSGN/n1749 ), .B(\UPIF/CSGN/n1752 ) );
    snl_nand02x1 \UPIF/CSGN/U1715  ( .ZN(\UPIF/CSGN/n1713 ), .A(ph_filewr_h), 
        .B(wacc) );
    snl_invx2 \UPIF/CSGN/U1557  ( .ZN(\pk_rread_h[41] ), .A(\UPIF/CSGN/n1695 )
         );
    snl_nor03x4 \UPIF/CSGN/U1570  ( .ZN(\pk_rread_h[0] ), .A(\UPIF/CSGN/n1649 
        ), .B(\UPIF/CSGN/n1648 ), .C(\UPIF/CSGN/n1653 ) );
    snl_nor02x1 \UPIF/CSGN/U1577  ( .ZN(pr_write_h), .A(\UPIF/CSGN/n1650 ), 
        .B(\UPIF/CSGN/n1652 ) );
    snl_nand03x0 \UPIF/CSGN/U1647  ( .ZN(\UPIF/CSGN/n1689 ), .A(
        \UPIF/CSGN/n1649 ), .B(\UPIF/CSGN/n1727 ), .C(\UPIF/CSGN/n1735 ) );
    snl_nand02x1 \UPIF/CSGN/U1660  ( .ZN(\UPIF/CSGN/n1663 ), .A(
        \UPIF/CSGN/n1743 ), .B(\UPIF/CSGN/n1737 ) );
    snl_and02x1 \UPIF/CSGN/U1640  ( .Z(\UPIF/CSGN/n1733 ), .A(
        \UPIF/CSGN/n1723 ), .B(\UPIF/CSGN/n1649 ) );
    snl_and02x1 \UPIF/CSGN/U1667  ( .Z(\UPIF/CSGN/n1747 ), .A(PA[7]), .B(
        \UPIF/CSGN/n1724 ) );
    snl_nor03x0 \UPIF/CSGN/U1609  ( .ZN(\pk_rwrit_h[18] ), .A(
        \UPIF/CSGN/n1696 ), .B(\UPIF/CSGN/n1665 ), .C(\UPIF/CSGN/n1639 ) );
    snl_nor02x1 \UPIF/CSGN/U1595  ( .ZN(\pk_rwrit_h[3] ), .A(\UPIF/CSGN/n1639 
        ), .B(\UPIF/CSGN/n1677 ) );
    snl_nand02x1 \UPIF/CSGN/U1682  ( .ZN(\UPIF/CSGN/n1710 ), .A(
        \UPIF/CSGN/n1750 ), .B(\UPIF/CSGN/n1728 ) );
    snl_nor03x0 \UPIF/CSGN/U1712  ( .ZN(\UPIF/CSGN/n1716 ), .A(PA[31]), .B(PA
        [26]), .C(PA[30]) );
    snl_nand02x1 \UPIF/CSGN/U1635  ( .ZN(\UPIF/CSGN/n1659 ), .A(
        \UPIF/CSGN/n1731 ), .B(\UPIF/CSGN/n1724 ) );
    snl_nand02x1 \UPIF/CSGN/U1699  ( .ZN(\UPIF/CSGN/n1705 ), .A(
        \UPIF/CSGN/n1756 ), .B(\UPIF/CSGN/n1732 ) );
    snl_invx05 \UPIF/CSGN/U1735  ( .ZN(\UPIF/CSGN/n1737 ), .A(
        \UPIF/CSGN/n1645 ) );
    snl_nor02x1 \UPIF/CSGN/U1709  ( .ZN(mem_cnfg_h), .A(\UPIF/CSGN/n1699 ), 
        .B(\UPIF/CSGN/n1679 ) );
    snl_nor02x3 \UPIF/CSGN/U1505  ( .ZN(\pk_rwrit_h[8] ), .A(\UPIF/CSGN/n1650 
        ), .B(\UPIF/CSGN/n1669 ) );
    snl_nor02x3 \UPIF/CSGN/U1522  ( .ZN(\pk_rread_h[9] ), .A(\UPIF/CSGN/n1664 
        ), .B(\UPIF/CSGN/n1654 ) );
    snl_nor02x1 \UPIF/CSGN/U1612  ( .ZN(\pk_rwrit_h[46] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1702 ) );
    snl_bufx1 \UPIF/CSGN/U1471  ( .Z(\UPIF/CSGN/n1638 ), .A(ad_latch) );
    snl_and02x2 \UPIF/CSGN/U1479  ( .Z(\pk_rread_h[39] ), .A(\UPIF/CSGN/n1745 
        ), .B(\UPIF/CSGN/n1743 ) );
    snl_and02x2 \UPIF/CSGN/U1487  ( .Z(\pk_rread_h[47] ), .A(PA[10]), .B(
        \UPIF/CSGN/reg_stat_h ) );
    snl_nor02x3 \UPIF/CSGN/U1517  ( .ZN(\pk_rread_h[16] ), .A(
        \UPIF/CSGN/n1671 ), .B(\UPIF/CSGN/n1700 ) );
    snl_nor02x1 \UPIF/CSGN/U1579  ( .ZN(ret_cont_wr), .A(\UPIF/CSGN/n1650 ), 
        .B(\UPIF/CSGN/n1659 ) );
    snl_nor02x1 \UPIF/CSGN/U1649  ( .ZN(\UPIF/CSGN/n1738 ), .A(
        \UPIF/CSGN/n1676 ), .B(PA[7]) );
    snl_nand02x1 \UPIF/CSGN/U1627  ( .ZN(\UPIF/CSGN/n1647 ), .A(PA[4]), .B(
        \UPIF/CSGN/n1728 ) );
    snl_invx1 \UPIF/CSGN/U1530  ( .ZN(seg_cnfg_h), .A(\UPIF/CSGN/n1658 ) );
    snl_invx2 \UPIF/CSGN/U1545  ( .ZN(\pk_rread_h[31] ), .A(\UPIF/CSGN/n1710 )
         );
    snl_invx2 \UPIF/CSGN/U1562  ( .ZN(\pk_rread_h[2] ), .A(\UPIF/CSGN/n1672 )
         );
    snl_nor03x0 \UPIF/CSGN/U1587  ( .ZN(\pk_rwrit_h[16] ), .A(
        \UPIF/CSGN/n1670 ), .B(\UPIF/CSGN/n1639 ), .C(\UPIF/CSGN/n1671 ) );
    snl_nor02x1 \UPIF/CSGN/U1600  ( .ZN(ph_ex2regwt_h), .A(\UPIF/CSGN/n1684 ), 
        .B(\UPIF/CSGN/n1685 ) );
    snl_nand02x1 \UPIF/CSGN/U1690  ( .ZN(\UPIF/CSGN/n1691 ), .A(
        \UPIF/CSGN/n1749 ), .B(\UPIF/CSGN/n1754 ) );
    snl_nand02x1 \UPIF/CSGN/U1700  ( .ZN(\UPIF/CSGN/n1682 ), .A(
        \UPIF/CSGN/n1755 ), .B(\UPIF/CSGN/n1753 ) );
    snl_invx05 \UPIF/CSGN/U1727  ( .ZN(\UPIF/CSGN/n1752 ), .A(
        \UPIF/CSGN/n1647 ) );
    snl_and02x1 \UPIF/CSGN/U1652  ( .Z(\UPIF/CSGN/n1740 ), .A(
        \UPIF/CSGN/n1739 ), .B(\UPIF/CSGN/n1649 ) );
    snl_nand02x1 \UPIF/CSGN/U1675  ( .ZN(\UPIF/CSGN/n1673 ), .A(
        \UPIF/CSGN/n1748 ), .B(\UPIF/CSGN/n1743 ) );
    snl_ao012x2 \UPIF/CSGN/U1476  ( .Z(\pk_rwrit_h[53] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[45] ), .C(ph_stregwt_h) );
    snl_and02x2 \UPIF/CSGN/U1478  ( .Z(\pk_rwrit_h[10] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[10] ) );
    snl_nor02x2 \UPIF/CSGN/U1494  ( .ZN(\pk_rwrit_h[34] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1667 ) );
    snl_nor02x3 \UPIF/CSGN/U1504  ( .ZN(\pk_rwrit_h[37] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1686 ) );
    snl_nor03x0 \UPIF/CSGN/U1634  ( .ZN(\UPIF/CSGN/n1731 ), .A(
        \UPIF/CSGN/n1648 ), .B(PA[6]), .C(\UPIF/CSGN/n1727 ) );
    snl_nand02x1 \UPIF/CSGN/U1698  ( .ZN(\UPIF/CSGN/n1674 ), .A(
        \UPIF/CSGN/n1756 ), .B(\UPIF/CSGN/n1724 ) );
    snl_nand02x1 \UPIF/CSGN/U1708  ( .ZN(\UPIF/CSGN/n1641 ), .A(
        \UPIF/CSGN/n1744 ), .B(\UPIF/CSGN/n1741 ) );
    snl_nor02x3 \UPIF/CSGN/U1523  ( .ZN(\pk_rread_h[10] ), .A(
        \UPIF/CSGN/n1696 ), .B(\UPIF/CSGN/n1654 ) );
    snl_invx2 \UPIF/CSGN/U1538  ( .ZN(\pk_rread_h[12] ), .A(\UPIF/CSGN/n1708 )
         );
    snl_nor02x1 \UPIF/CSGN/U1608  ( .ZN(\pk_rwrit_h[49] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1695 ) );
    snl_and02x1 \UPIF/CSGN/U1613  ( .Z(\pk_rwrit_h[23] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[16] ) );
    snl_invx2 \UPIF/CSGN/U1544  ( .ZN(\pk_rread_h[35] ), .A(\UPIF/CSGN/n1673 )
         );
    snl_invx2 \UPIF/CSGN/U1556  ( .ZN(\pk_rread_h[25] ), .A(\UPIF/CSGN/n1691 )
         );
    snl_invx2 \UPIF/CSGN/U1571  ( .ZN(\pk_rread_h[55] ), .A(\UPIF/CSGN/n1663 )
         );
    snl_nor03x0 \UPIF/CSGN/U1594  ( .ZN(\pk_rwrit_h[15] ), .A(
        \UPIF/CSGN/n1670 ), .B(\UPIF/CSGN/n1676 ), .C(\UPIF/CSGN/n1639 ) );
    snl_nand02x1 \UPIF/CSGN/U1683  ( .ZN(\UPIF/CSGN/n1653 ), .A(
        \UPIF/CSGN/n1734 ), .B(PA[4]) );
    snl_nor04x0 \UPIF/CSGN/U1713  ( .ZN(\UPIF/CSGN/n1759 ), .A(PA[20]), .B(PA
        [21]), .C(PA[28]), .D(\UPIF/CSGN/n1644 ) );
    snl_invx05 \UPIF/CSGN/U1734  ( .ZN(\UPIF/CSGN/n1745 ), .A(
        \UPIF/CSGN/n1688 ) );
    snl_nand12x1 \UPIF/CSGN/U1641  ( .ZN(\UPIF/CSGN/n1671 ), .A(PA[3]), .B(
        \UPIF/CSGN/n1726 ) );
    snl_nand02x1 \UPIF/CSGN/U1666  ( .ZN(\UPIF/CSGN/n1688 ), .A(
        \UPIF/CSGN/n1734 ), .B(PA[7]) );
    snl_invx2 \UPIF/CSGN/U1563  ( .ZN(\pk_rread_h[34] ), .A(\UPIF/CSGN/n1655 )
         );
    snl_and02x1 \UPIF/CSGN/U1653  ( .Z(\UPIF/CSGN/n1741 ), .A(
        \UPIF/CSGN/n1724 ), .B(\UPIF/CSGN/n1722 ) );
    snl_nand02x1 \UPIF/CSGN/U1674  ( .ZN(\UPIF/CSGN/n1706 ), .A(
        \UPIF/CSGN/n1747 ), .B(\UPIF/CSGN/n1743 ) );
    snl_nor02x2 \UPIF/CSGN/U1481  ( .ZN(\pk_rwrit_h[33] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1661 ) );
    snl_and02x2 \UPIF/CSGN/U1486  ( .Z(\pk_rread_h[60] ), .A(\UPIF/CSGN/n1740 
        ), .B(\UPIF/CSGN/n1738 ) );
    snl_nor02x1 \UPIF/CSGN/U1586  ( .ZN(\pk_rwrit_h[64] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1666 ) );
    snl_and23x0 \UPIF/CSGN/U1691  ( .Z(\UPIF/CSGN/n1755 ), .A(
        \UPIF/CSGN/n1649 ), .B(PA[7]), .C(\UPIF/CSGN/n1729 ) );
    snl_nand02x1 \UPIF/CSGN/U1701  ( .ZN(\UPIF/CSGN/n1693 ), .A(
        \UPIF/CSGN/n1755 ), .B(\UPIF/CSGN/n1754 ) );
    snl_invx05 \UPIF/CSGN/U1626  ( .ZN(\UPIF/CSGN/n1727 ), .A(PA[4]) );
    snl_invx05 \UPIF/CSGN/U1726  ( .ZN(\UPIF/CSGN/n1744 ), .A(
        \UPIF/CSGN/n1646 ) );
    snl_nor02x3 \UPIF/CSGN/U1511  ( .ZN(seg_config_wr), .A(\UPIF/CSGN/n1650 ), 
        .B(\UPIF/CSGN/n1658 ) );
    snl_nor02x3 \UPIF/CSGN/U1516  ( .ZN(\pk_rread_h[53] ), .A(
        \UPIF/CSGN/n1645 ), .B(\UPIF/CSGN/n1646 ) );
    snl_ao1b1b3x2 \UPIF/CSGN/U1531  ( .Z(\pk_rwrit_h[50] ), .A(
        \UPIF/CSGN/n1711 ), .B(phsaerrh), .C(ph_dregsl_h), .D(
        \UPIF/CSGN/n1712 ), .E(ph_stdatlth) );
    snl_invx2 \UPIF/CSGN/U1536  ( .ZN(\pk_rread_h[40] ), .A(\UPIF/CSGN/n1701 )
         );
    snl_invx2 \UPIF/CSGN/U1558  ( .ZN(\pk_rread_h[33] ), .A(\UPIF/CSGN/n1668 )
         );
    snl_nor03x0 \UPIF/CSGN/U1578  ( .ZN(\pk_rwrit_h[14] ), .A(
        \UPIF/CSGN/n1653 ), .B(\UPIF/CSGN/n1639 ), .C(\UPIF/CSGN/n1654 ) );
    snl_nor03x0 \UPIF/CSGN/U1601  ( .ZN(\UPIF/CSGN/n_1047 ), .A(
        \UPIF/CSGN/n1641 ), .B(WR), .C(\UPIF/CSGN/n1642 ) );
    snl_nand02x1 \UPIF/CSGN/U1648  ( .ZN(\UPIF/CSGN/n1714 ), .A(
        \UPIF/CSGN/n1736 ), .B(\UPIF/CSGN/n1737 ) );
    snl_invx05 \UPIF/CSGN/U1668  ( .ZN(\UPIF/CSGN/n1711 ), .A(ph_srdalth) );
    snl_and02x1 \UPIF/CSGN/U1606  ( .Z(\pk_rwrit_h[45] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[37] ) );
    snl_and02x2 \UPIF/CSGN/U1488  ( .Z(\pk_rread_h[54] ), .A(\UPIF/CSGN/n1743 
        ), .B(\UPIF/CSGN/n1738 ) );
    snl_invx2 \UPIF/CSGN/U1543  ( .ZN(\pk_rread_h[32] ), .A(\UPIF/CSGN/n1660 )
         );
    snl_nor02x1 \UPIF/CSGN/U1581  ( .ZN(\pk_rwrit_h[63] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1662 ) );
    snl_nor02x1 \UPIF/CSGN/U1621  ( .ZN(\UPIF/CSGN/n1723 ), .A(
        \UPIF/CSGN/n1648 ), .B(PA[4]) );
    snl_nand02x1 \UPIF/CSGN/U1721  ( .ZN(\UPIF/CSGN/n1680 ), .A(
        \pk_rread_h[54] ), .B(\UPIF/reg_wr ) );
    snl_nand02x1 \UPIF/CSGN/U1696  ( .ZN(\UPIF/CSGN/n1707 ), .A(
        \UPIF/CSGN/n1755 ), .B(\UPIF/CSGN/n1751 ) );
    snl_nand02x1 \UPIF/CSGN/U1706  ( .ZN(\UPIF/CSGN/n1685 ), .A(
        \UPIF/CSGN/n1744 ), .B(\UPIF/CSGN/n1742 ) );
    snl_invx2 \UPIF/CSGN/U1551  ( .ZN(\pk_rread_h[51] ), .A(\UPIF/CSGN/n1692 )
         );
    snl_invx2 \UPIF/CSGN/U1564  ( .ZN(\pk_rread_h[6] ), .A(\UPIF/CSGN/n1690 )
         );
    snl_nand02x1 \UPIF/CSGN/U1654  ( .ZN(\UPIF/CSGN/n1666 ), .A(
        \UPIF/CSGN/n1741 ), .B(\UPIF/CSGN/n1736 ) );
    snl_nand02x1 \UPIF/CSGN/U1673  ( .ZN(\UPIF/CSGN/n1702 ), .A(
        \UPIF/CSGN/n1746 ), .B(\UPIF/CSGN/n1743 ) );
    snl_nor02x1 \UPIF/CSGN/U1576  ( .ZN(\pk_rwrit_h[61] ), .A(
        \UPIF/CSGN/n1639 ), .B(\UPIF/CSGN/n1651 ) );
    snl_nand02x1 \UPIF/CSGN/U1646  ( .ZN(\UPIF/CSGN/n1645 ), .A(
        \UPIF/CSGN/n1734 ), .B(\UPIF/CSGN/n1722 ) );
    snl_nand02x1 \UPIF/CSGN/U1661  ( .ZN(\UPIF/CSGN/n1687 ), .A(
        \UPIF/CSGN/n1731 ), .B(\UPIF/CSGN/n1728 ) );
    snl_invx05 \UPIF/CSGN/U1628  ( .ZN(\UPIF/CSGN/n1721 ), .A(PA[8]) );
    snl_nor02x2 \UPIF/CSGN/U1493  ( .ZN(\pk_rwrit_h[25] ), .A(
        \UPIF/CSGN/n1650 ), .B(\UPIF/CSGN/n1682 ) );
    snl_nor02x3 \UPIF/CSGN/U1518  ( .ZN(\pk_rread_h[15] ), .A(
        \UPIF/CSGN/n1700 ), .B(\UPIF/CSGN/n1676 ) );
    snl_nor02x3 \UPIF/CSGN/U1524  ( .ZN(\pk_rread_h[14] ), .A(
        \UPIF/CSGN/n1653 ), .B(\UPIF/CSGN/n1665 ) );
    snl_and02x1 \UPIF/CSGN/U1588  ( .Z(\pk_rwrit_h[22] ), .A(\UPIF/reg_wr ), 
        .B(\pk_rread_h[15] ) );
    snl_and02x1 \UPIF/CSGN/U1593  ( .Z(cnfg_write_h), .A(\UPIF/reg_wr ), .B(
        mem_cnfg_h) );
    snl_invx05 \UPIF/CSGN/U1733  ( .ZN(\UPIF/CSGN/n1746 ), .A(
        \UPIF/CSGN/n1683 ) );
    snl_nand02x1 \UPIF/CSGN/U1684  ( .ZN(\UPIF/CSGN/n1686 ), .A(
        \UPIF/CSGN/n1751 ), .B(\UPIF/CSGN/n1749 ) );
    snl_nand04x0 \UPIF/CSGN/U1714  ( .ZN(\UPIF/CSGN/n1719 ), .A(PA[27]), .B(PA
        [29]), .C(PA[13]), .D(\UPIF/CSGN/n1759 ) );
    snl_ao023x1 \UPIF/CSGN/U1614  ( .Z(\pk_rwrit_h[67] ), .A(ph_filewr_h), .B(
        \UPIF/CSGN/n1704 ), .C(wexacc), .D(\pk_rread_h[62] ), .E(\UPIF/reg_wr 
        ) );
    snl_invx05 \UPIF/CSGN/U1728  ( .ZN(\UPIF/CSGN/n1751 ), .A(
        \UPIF/CSGN/n1653 ) );
    snl_nor02x3 \UPIF/CSGN/U1503  ( .ZN(\pk_rwrit_h[6] ), .A(\UPIF/CSGN/n1650 
        ), .B(\UPIF/CSGN/n1690 ) );
    snl_nand02x1 \UPIF/CSGN/U1633  ( .ZN(\UPIF/CSGN/n1658 ), .A(
        \UPIF/CSGN/n1730 ), .B(\UPIF/CSGN/n1724 ) );
    snl_and02x1 \LBUS/ldoecnt_5/U8  ( .Z(ph_ldaoutenhp), .A(ph_lbwrh), .B(
        \LBUS/temp[3] ) );
    snl_mux21x1 \ADOSEL/seladr_2/U10  ( .Z(LOUT[15]), .A(\pgsadrh[15] ), .B(
        \pgmuxout[15] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U12  ( .Z(LOUT[13]), .A(\pgsadrh[13] ), .B(
        \pgmuxout[13] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U13  ( .Z(LOUT[12]), .A(\pgsadrh[12] ), .B(
        \pgmuxout[12] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U14  ( .Z(LOUT[11]), .A(\pgsadrh[11] ), .B(
        \pgmuxout[11] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U15  ( .Z(LOUT[10]), .A(\pgsadrh[10] ), .B(
        \pgmuxout[10] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U17  ( .Z(LOUT[8]), .A(\pgsadrh[8] ), .B(
        \pgmuxout[8] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U11  ( .Z(LOUT[14]), .A(\pgsadrh[14] ), .B(
        \pgmuxout[14] ), .S(ph_ldaoutenh2) );
    snl_mux21x1 \ADOSEL/seladr_2/U16  ( .Z(LOUT[9]), .A(\pgsadrh[9] ), .B(
        \pgmuxout[9] ), .S(ph_ldaoutenh2) );
    snl_and02x1 \CONS/phinc20_1/U6  ( .Z(\CONS/phinc20_1/gg_out[3] ), .A(
        \CONS/phinc20_1/gp_out[3] ), .B(\CONS/phinc20_1/gg_out[2] ) );
    snl_and02x1 \CONS/phinc20_1/U7  ( .Z(\CONS/phinc20_1/gg_out[1] ), .A(
        \CONS/phinc20_1/gp_out[1] ), .B(\CONS/phinc20_1/gp_out[0] ) );
    snl_and02x1 \CONS/phinc20_1/U8  ( .Z(\CONS/phinc20_1/gg_out[2] ), .A(
        \CONS/phinc20_1/gp_out[2] ), .B(\CONS/phinc20_1/gg_out[1] ) );
    snl_and02x1 \CODEIF/inc19_1/U6  ( .Z(\CODEIF/pgctrinc[15] ), .A(
        \CODEIF/inc19_1/n3763 ), .B(\CODEIF/inc19_1/n3764 ) );
    snl_and02x1 \CODEIF/inc19_1/U7  ( .Z(\CODEIF/inc19_1/gg_out[3] ), .A(
        \CODEIF/inc19_1/gp_out[3] ), .B(\CODEIF/inc19_1/gg_out[2] ) );
    snl_and02x1 \CODEIF/inc19_1/U8  ( .Z(\CODEIF/inc19_1/gg_out[1] ), .A(
        \CODEIF/inc19_1/gp_out[1] ), .B(\CODEIF/inc19_1/gp_out[0] ) );
    snl_and02x1 \CODEIF/inc19_1/U9  ( .Z(\CODEIF/inc19_1/gg_out[2] ), .A(
        \CODEIF/inc19_1/gp_out[2] ), .B(\CODEIF/inc19_1/gg_out[1] ) );
    snl_and02x1 \LBUS/ldoecnt_2/U8  ( .Z(ph_ldaoutenh2), .A(ph_lbwrh), .B(
        \LBUS/temp[3] ) );
    snl_and02x1 \UPIF/RCTL/U121  ( .Z(pol_status), .A(\UPIF/RCTL/n1031 ), .B(
        \UPIF/RCTL/n1023 ) );
    snl_nor02x1 \UPIF/RCTL/U126  ( .ZN(\UPIF/RCTL/n1034 ), .A(
        \UPIF/RCTL/irt[1] ), .B(\UPIF/RCTL/irt[0] ) );
    snl_invx05 \UPIF/RCTL/U134  ( .ZN(\UPIF/RCTL/n1033 ), .A(
        \UPIF/RCTL/irt[1] ) );
    snl_nand13x1 \UPIF/RCTL/U141  ( .ZN(\UPIF/RCTL/n1041 ), .A(PA[12]), .B(PA
        [11]), .C(PA[13]) );
    snl_invx05 \UPIF/RCTL/U148  ( .ZN(\UPIF/RCTL/nrt[1] ), .A(
        \UPIF/RCTL/n1027 ) );
    snl_nor08x1 \UPIF/RCTL/U114  ( .ZN(\UPIF/RCTL/n1023 ), .A(PA[26]), .B(PA
        [25]), .C(PA[24]), .D(PA[31]), .E(PA[30]), .F(PA[28]), .G(
        \UPIF/RCTL/n1037 ), .H(\UPIF/RCTL/n1038 ) );
    snl_oa013x1 \UPIF/RCTL/U128  ( .Z(\UPIF/ph_accessenh ), .A(
        \UPIF/RCTL/irt[2] ), .B(\UPIF/RCTL/irt[3] ), .C(\UPIF/RCTL/n_831 ), 
        .D(\UPIF/RCTL/reg_file_h ) );
    snl_nor03x0 \UPIF/RCTL/U133  ( .ZN(\UPIF/RCTL/*cell*4328/U25/CONTROL2 ), 
        .A(\UPIF/RCTL/irt[2] ), .B(\UPIF/RCTL/irt[1] ), .C(\UPIF/RCTL/n1036 )
         );
    snl_oa113x1 \UPIF/RCTL/U146  ( .Z(\UPIF/RCTL/n1042 ), .A(code_area_h), .B(
        \UPIF/RCTL/n1023 ), .C(\UPIF/RCTL/reg_file_h ), .D(\UPIF/RCTL/n1034 ), 
        .E(ADS) );
    snl_nor02x2 \UPIF/RCTL/U115  ( .ZN(cif_cont), .A(\UPIF/RCTL/n1025 ), .B(
        \UPIF/RCTL/n1032 ) );
    snl_ao022x1 \UPIF/RCTL/U120  ( .Z(\UPIF/RCTL/reg_eoc ), .A(
        \UPIF/RCTL/irt[0] ), .B(\UPIF/RCTL/irt[1] ), .C(\UPIF/RCTL/irt[2] ), 
        .D(\UPIF/iready ) );
    snl_invx05 \UPIF/RCTL/U132  ( .ZN(\UPIF/RCTL/n1036 ), .A(
        \UPIF/RCTL/irt[0] ) );
    snl_oai122x0 \UPIF/RCTL/U116  ( .ZN(\UPIF/RCTL/nrt[0] ), .A(IBSY), .B(
        \UPIF/RCTL/n1024 ), .C(\UPIF/iready ), .D(\UPIF/RCTL/n1025 ), .E(
        \UPIF/RCTL/n1026 ) );
    snl_aoi012x1 \UPIF/RCTL/U117  ( .ZN(\UPIF/RCTL/n1027 ), .A(
        \UPIF/RCTL/n1025 ), .B(\UPIF/RCTL/irt[0] ), .C(\UPIF/RCTL/reg_eoc ) );
    snl_nor02x1 \UPIF/RCTL/U119  ( .ZN(\UPIF/RCTL/nrt[3] ), .A(
        \UPIF/RCTL/n1024 ), .B(\UPIF/RCTL/n1030 ) );
    snl_nand12x1 \UPIF/RCTL/U127  ( .ZN(\UPIF/RCTL/n_839 ), .A(
        \UPIF/RCTL/nrt[0] ), .B(\UPIF/RCTL/n1027 ) );
    snl_oai122x0 \UPIF/RCTL/U129  ( .ZN(\UPIF/RCTL/n1031 ), .A(
        \UPIF/RCTL/n1033 ), .B(\UPIF/RCTL/irt[0] ), .C(\UPIF/RCTL/n1035 ), .D(
        IBSY), .E(\UPIF/RCTL/n1025 ) );
    snl_nor02x1 \UPIF/RCTL/U147  ( .ZN(\UPIF/RCTL/n1024 ), .A(
        \UPIF/RCTL/irt[3] ), .B(\UPIF/RCTL/n1042 ) );
    snl_ffqrnx1 \UPIF/RCTL/irt_reg[1]  ( .Q(\UPIF/RCTL/irt[1] ), .D(
        \UPIF/RCTL/nrt[1] ), .RN(n10733), .CP(SCLK) );
    snl_invx05 \UPIF/RCTL/U135  ( .ZN(\UPIF/RCTL/n1025 ), .A(
        \UPIF/RCTL/irt[2] ) );
    snl_and34x0 \UPIF/RCTL/U140  ( .Z(\UPIF/RCTL/n1040 ), .A(PA[15]), .B(PA
        [14]), .C(PA[16]), .D(\UPIF/RCTL/n1039 ) );
    snl_ffqrnx1 \UPIF/RCTL/irt_reg[3]  ( .Q(\UPIF/RCTL/irt[3] ), .D(
        \UPIF/RCTL/nrt[3] ), .RN(n10733), .CP(SCLK) );
    snl_sffqrnx1 \UPIF/RCTL/reg_wr_reg  ( .Q(\UPIF/reg_wr ), .D(1'b0), .RN(
        n10733), .SD(\UPIF/RCTL/*cell*4328/U25/CONTROL2 ), .SE(WR), .CP(SCLK)
         );
    snl_invx05 \UPIF/RCTL/U137  ( .ZN(\UPIF/RCTL/n1030 ), .A(IBSY) );
    snl_nand14x0 \UPIF/RCTL/U142  ( .ZN(\UPIF/RCTL/n1038 ), .A(
        \UPIF/RCTL/n1041 ), .B(PA[27]), .C(PA[29]), .D(\UPIF/RCTL/n1040 ) );
    snl_sffqqnrnx1 \UPIF/RCTL/rdy_oe_h_reg  ( .QN(RDYOLCNT), .D(
        \UPIF/RCTL/n_831 ), .RN(n10733), .SD(1'b1), .SE(\UPIF/RCTL/irt[2] ), 
        .CP(SCLK) );
    snl_and02x1 \UPIF/RCTL/U122  ( .Z(cif_byte), .A(\UPIF/RCTL/irt[2] ), .B(
        \UPIF/write_by_h ) );
    snl_invx05 \UPIF/RCTL/U125  ( .ZN(\UPIF/RCTL/n_837 ), .A(WR) );
    snl_ffqrnx1 \UPIF/RCTL/irt_reg[2]  ( .Q(\UPIF/RCTL/irt[2] ), .D(
        \UPIF/RCTL/nrt[2] ), .RN(n10733), .CP(SCLK) );
    snl_sffqqnrnx1 \UPIF/RCTL/pdoe_reg  ( .QN(PDCNT), .D(1'b0), .RN(n10733), 
        .SD(\UPIF/RCTL/n_839 ), .SE(\UPIF/RCTL/n_837 ), .CP(SCLK) );
    snl_nor02x1 \UPIF/RCTL/U139  ( .ZN(\UPIF/RCTL/n1039 ), .A(PA[18]), .B(PA
        [17]) );
    snl_ffqrnx1 \UPIF/RCTL/irt_reg[0]  ( .Q(\UPIF/RCTL/irt[0] ), .D(
        \UPIF/RCTL/nrt[0] ), .RN(n10733), .CP(SCLK) );
    snl_ffqrnx1 \UPIF/RCTL/ready_eoc_reg  ( .Q(\UPIF/ready_eoc ), .D(
        \UPIF/RCTL/reg_eoc ), .RN(n10733), .CP(SCLK) );
    snl_invx05 \UPIF/RCTL/U145  ( .ZN(\UPIF/RCTL/n_831 ), .A(\UPIF/RCTL/n1034 
        ) );
    snl_nor02x1 \UPIF/RCTL/U123  ( .ZN(\UPIF/tr_count_lt ), .A(WR), .B(
        \UPIF/RCTL/n1026 ) );
    snl_aoi113x0 \UPIF/RCTL/U130  ( .ZN(\UPIF/RCTL/n1029 ), .A(
        \UPIF/RCTL/reg_file_h ), .B(WR), .C(\UPIF/write_by_h ), .D(
        \UPIF/RCTL/n1023 ), .E(code_area_h) );
    snl_or05x1 \UPIF/RCTL/U138  ( .Z(\UPIF/RCTL/n1037 ), .A(PA[23]), .B(PA[22]
        ), .C(PA[21]), .D(PA[20]), .E(PA[19]) );
    snl_ffqnrnx2 \UPIF/RCTL/ready_cpu_reg  ( .QN(RDYOL), .D(
        \UPIF/RCTL/reg_eoc ), .RN(n10733), .CP(SCLK) );
    snl_oai023x0 \UPIF/RCTL/U118  ( .ZN(\UPIF/RCTL/nrt[2] ), .A(
        \UPIF/RCTL/n1028 ), .B(IBSY), .C(\UPIF/RCTL/n1029 ), .D(\UPIF/iready ), 
        .E(\UPIF/RCTL/n1025 ) );
    snl_nor03x0 \UPIF/RCTL/U124  ( .ZN(ph_cperlt_h), .A(\UPIF/RCTL/n1032 ), 
        .B(\UPIF/RCTL/irt[0] ), .C(\UPIF/RCTL/n1033 ) );
    snl_aoi012x1 \UPIF/RCTL/U131  ( .ZN(\UPIF/RCTL/n1028 ), .A(ADS), .B(
        \UPIF/RCTL/n1034 ), .C(\UPIF/RCTL/irt[3] ) );
    snl_invx05 \UPIF/RCTL/U136  ( .ZN(\UPIF/RCTL/n1032 ), .A(code_area_h) );
    snl_invx05 \UPIF/RCTL/U143  ( .ZN(\UPIF/RCTL/n1026 ), .A(
        \UPIF/RCTL/*cell*4328/U25/CONTROL2 ) );
    snl_aoi012x1 \UPIF/RCTL/U144  ( .ZN(\UPIF/RCTL/n1035 ), .A(
        \UPIF/RCTL/n1036 ), .B(ADS), .C(\UPIF/RCTL/irt[3] ) );
    snl_aoi023x0 \CONS/lte_124/U6  ( .ZN(\CONS/n300 ), .A(\CONS/lte_124/n63 ), 
        .B(\CONS/lte_124/n64 ), .C(\CONS/lte_124/n65 ), .D(\pk_pc_h[18] ), .E(
        \CONS/lte_124/n66 ) );
    snl_and02x1 \CONS/lte_124/U14  ( .Z(\CONS/lte_124/n293 ), .A(
        \CONS/lte_124/n294 ), .B(\pk_pcs2_h[12] ) );
    snl_invx05 \CONS/lte_124/U21  ( .ZN(\CONS/lte_124/n68 ), .A(\pk_pcs2_h[3] 
        ) );
    snl_invx05 \CONS/lte_124/U28  ( .ZN(\CONS/lte_124/n292 ), .A(
        \pk_pcs2_h[10] ) );
    snl_invx05 \CONS/lte_124/U33  ( .ZN(\CONS/lte_124/n300 ), .A(
        \pk_pcs2_h[15] ) );
    snl_aoi22b2x0 \CONS/lte_124/U7  ( .ZN(\CONS/lte_124/n67 ), .A(
        \CONS/lte_124/n70 ), .B(\pk_pcs2_h[2] ), .C(\pk_pc_h[3] ), .D(
        \CONS/lte_124/n68 ), .E(\pk_pc_h[2] ), .F(\CONS/lte_124/n69 ) );
    snl_and02x1 \CONS/lte_124/U8  ( .Z(\CONS/lte_124/n71 ), .A(
        \CONS/lte_124/n72 ), .B(\pk_pcs2_h[4] ) );
    snl_aoi223x0 \CONS/lte_124/U13  ( .ZN(\CONS/lte_124/n287 ), .A(
        \CONS/lte_124/n288 ), .B(\CONS/lte_124/n289 ), .C(\CONS/lte_124/n290 ), 
        .D(\pk_pc_h[11] ), .E(\CONS/lte_124/n291 ), .F(\pk_pc_h[10] ), .G(
        \CONS/lte_124/n292 ) );
    snl_invx05 \CONS/lte_124/U34  ( .ZN(\CONS/lte_124/n303 ), .A(\pk_pc_h[16] 
        ) );
    snl_nand02x1 \CONS/lte_124/U41  ( .ZN(\CONS/lte_124/n281 ), .A(
        \pk_pcs2_h[5] ), .B(\CONS/lte_124/n307 ) );
    snl_nand12x1 \CONS/lte_124/U46  ( .ZN(\CONS/lte_124/n297 ), .A(
        \pk_pc_h[14] ), .B(\pk_pcs2_h[14] ) );
    snl_invx05 \CONS/lte_124/U26  ( .ZN(\CONS/lte_124/n285 ), .A(\pk_pc_h[8] )
         );
    snl_oai223x0 \CONS/lte_124/U48  ( .ZN(\CONS/lte_124/n64 ), .A(
        \CONS/lte_124/n304 ), .B(\CONS/lte_124/n296 ), .C(\CONS/lte_124/n302 ), 
        .D(\pk_pcs2_h[16] ), .E(\CONS/lte_124/n303 ), .F(\pk_pcs2_h[17] ), .G(
        \CONS/lte_124/n310 ) );
    snl_nor02x1 \CONS/lte_124/U9  ( .ZN(\CONS/lte_124/n73 ), .A(\pk_pc_h[3] ), 
        .B(\CONS/lte_124/n68 ) );
    snl_nor02x1 \CONS/lte_124/U12  ( .ZN(\CONS/lte_124/n286 ), .A(\pk_pc_h[7] 
        ), .B(\CONS/lte_124/n282 ) );
    snl_invx05 \CONS/lte_124/U35  ( .ZN(\CONS/lte_124/n310 ), .A(\pk_pc_h[17] 
        ) );
    snl_invx05 \CONS/lte_124/U27  ( .ZN(\CONS/lte_124/n308 ), .A(\pk_pc_h[9] )
         );
    snl_nand12x1 \CONS/lte_124/U40  ( .ZN(\CONS/lte_124/n279 ), .A(
        \pk_pc_h[6] ), .B(\pk_pcs2_h[6] ) );
    snl_aoi022x1 \CONS/lte_124/U20  ( .ZN(\CONS/lte_124/n70 ), .A(\pk_pc_h[1] 
        ), .B(\CONS/lte_124/n305 ), .C(\CONS/lte_124/n306 ), .D(\pk_pc_h[0] )
         );
    snl_nand12x1 \CONS/lte_124/U49  ( .ZN(\CONS/lte_124/n63 ), .A(
        \pk_pc_h[18] ), .B(\pk_pcs2_h[18] ) );
    snl_invx05 \CONS/lte_124/U29  ( .ZN(\CONS/lte_124/n291 ), .A(
        \pk_pcs2_h[11] ) );
    snl_nand02x1 \CONS/lte_124/U47  ( .ZN(\CONS/lte_124/n299 ), .A(
        \pk_pcs2_h[13] ), .B(\CONS/lte_124/n309 ) );
    snl_aoi223x0 \CONS/lte_124/U10  ( .ZN(\CONS/lte_124/n278 ), .A(
        \CONS/lte_124/n279 ), .B(\CONS/lte_124/n280 ), .C(\CONS/lte_124/n281 ), 
        .D(\pk_pc_h[7] ), .E(\CONS/lte_124/n282 ), .F(\pk_pc_h[6] ), .G(
        \CONS/lte_124/n283 ) );
    snl_nor02x1 \CONS/lte_124/U15  ( .ZN(\CONS/lte_124/n295 ), .A(
        \pk_pc_h[11] ), .B(\CONS/lte_124/n291 ) );
    snl_and02x1 \CONS/lte_124/U17  ( .Z(\CONS/lte_124/n302 ), .A(
        \CONS/lte_124/n303 ), .B(\pk_pcs2_h[16] ) );
    snl_invx05 \CONS/lte_124/U22  ( .ZN(\CONS/lte_124/n72 ), .A(\pk_pc_h[4] )
         );
    snl_invx05 \CONS/lte_124/U32  ( .ZN(\CONS/lte_124/n301 ), .A(
        \pk_pcs2_h[14] ) );
    snl_oai223x0 \CONS/lte_124/U39  ( .ZN(\CONS/lte_124/n280 ), .A(
        \CONS/lte_124/n73 ), .B(\CONS/lte_124/n67 ), .C(\CONS/lte_124/n71 ), 
        .D(\pk_pcs2_h[4] ), .E(\CONS/lte_124/n72 ), .F(\pk_pcs2_h[5] ), .G(
        \CONS/lte_124/n307 ) );
    snl_invx05 \CONS/lte_124/U30  ( .ZN(\CONS/lte_124/n294 ), .A(\pk_pc_h[12] 
        ) );
    snl_oai223x0 \CONS/lte_124/U42  ( .ZN(\CONS/lte_124/n289 ), .A(
        \CONS/lte_124/n286 ), .B(\CONS/lte_124/n278 ), .C(\CONS/lte_124/n284 ), 
        .D(\pk_pcs2_h[8] ), .E(\CONS/lte_124/n285 ), .F(\pk_pcs2_h[9] ), .G(
        \CONS/lte_124/n308 ) );
    snl_oai223x0 \CONS/lte_124/U45  ( .ZN(\CONS/lte_124/n298 ), .A(
        \CONS/lte_124/n295 ), .B(\CONS/lte_124/n287 ), .C(\CONS/lte_124/n293 ), 
        .D(\pk_pcs2_h[12] ), .E(\CONS/lte_124/n294 ), .F(\pk_pcs2_h[13] ), .G(
        \CONS/lte_124/n309 ) );
    snl_and02x1 \CONS/lte_124/U11  ( .Z(\CONS/lte_124/n284 ), .A(
        \CONS/lte_124/n285 ), .B(\pk_pcs2_h[8] ) );
    snl_invx05 \CONS/lte_124/U19  ( .ZN(\CONS/lte_124/n305 ), .A(
        \pk_pcs2_h[1] ) );
    snl_invx05 \CONS/lte_124/U25  ( .ZN(\CONS/lte_124/n282 ), .A(
        \pk_pcs2_h[7] ) );
    snl_aoi01b2x1 \CONS/lte_124/U37  ( .ZN(\CONS/lte_124/n306 ), .A(
        \CONS/lte_124/n305 ), .B(\pk_pc_h[1] ), .C(\pk_pcs2_h[0] ) );
    snl_nand02x1 \CONS/lte_124/U50  ( .ZN(\CONS/lte_124/n65 ), .A(
        \pk_pcs2_h[17] ), .B(\CONS/lte_124/n310 ) );
    snl_aoi223x0 \CONS/lte_124/U16  ( .ZN(\CONS/lte_124/n296 ), .A(
        \CONS/lte_124/n297 ), .B(\CONS/lte_124/n298 ), .C(\CONS/lte_124/n299 ), 
        .D(\pk_pc_h[15] ), .E(\CONS/lte_124/n300 ), .F(\pk_pc_h[14] ), .G(
        \CONS/lte_124/n301 ) );
    snl_nor02x1 \CONS/lte_124/U18  ( .ZN(\CONS/lte_124/n304 ), .A(
        \pk_pc_h[15] ), .B(\CONS/lte_124/n300 ) );
    snl_invx05 \CONS/lte_124/U36  ( .ZN(\CONS/lte_124/n66 ), .A(
        \pk_pcs2_h[18] ) );
    snl_nand12x1 \CONS/lte_124/U43  ( .ZN(\CONS/lte_124/n288 ), .A(
        \pk_pc_h[10] ), .B(\pk_pcs2_h[10] ) );
    snl_invx05 \CONS/lte_124/U23  ( .ZN(\CONS/lte_124/n307 ), .A(\pk_pc_h[5] )
         );
    snl_invx05 \CONS/lte_124/U24  ( .ZN(\CONS/lte_124/n283 ), .A(
        \pk_pcs2_h[6] ) );
    snl_invx05 \CONS/lte_124/U31  ( .ZN(\CONS/lte_124/n309 ), .A(\pk_pc_h[13] 
        ) );
    snl_nand02x1 \CONS/lte_124/U38  ( .ZN(\CONS/lte_124/n69 ), .A(
        \pk_pcs2_h[2] ), .B(\CONS/lte_124/n70 ) );
    snl_nand02x1 \CONS/lte_124/U44  ( .ZN(\CONS/lte_124/n290 ), .A(
        \pk_pcs2_h[9] ), .B(\CONS/lte_124/n308 ) );
    snl_invx05 \SADR/ADRFF/U149  ( .ZN(\SADR/ADRFF/n9119 ), .A(n10732) );
    snl_invx1 \SADR/ADRFF/U153  ( .ZN(\SADR/ADRFF/n9123 ), .A(
        \SADR/ADRFF/n9122 ) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[27]  ( .Q(\pgsadrh[27] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[27] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[14]  ( .Q(\pgsadrh[14] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[14] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[2]  ( .Q(\pgsadrh[2] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprlh[5] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[6]  ( .Q(\SADR/m_fadrl[6] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[6] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[23]  ( .Q(\pgsadrh[23] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[23] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[10]  ( .Q(\pgsadrh[10] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[10] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[6]  ( .Q(\pgsadrh[6] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprlh[9] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_invx1 \SADR/ADRFF/U154  ( .ZN(\SADR/ADRFF/n9124 ), .A(
        \SADR/ADRFF/n9122 ) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[19]  ( .Q(\pgsadrh[19] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[19] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[25]  ( .Q(\pgsadrh[25] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[25] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[21]  ( .Q(\pgsadrh[21] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[21] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[12]  ( .Q(\pgsadrh[12] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[12] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[16]  ( .Q(\pgsadrh[16] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[16] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[9]  ( .Q(\pgsadrh[9] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgsdprlh[12] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[4]  ( .Q(\pgsadrh[4] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprlh[7] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[9]  ( .Q(\SADR/m_fadrl[9] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[9] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[0]  ( .Q(\pgsadrh[0] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[0] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[4]  ( .Q(\SADR/m_fadrl[4] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[4] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgbitnoh_reg[2]  ( .Q(\pgbitnoh[2] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/intbitno[2] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrh_reg[30]  ( .Q(\SADR/m_fadrh[30] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprhh[30] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrh_reg[29]  ( .Q(\SADR/m_fadrh[29] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprhh[29] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[22]  ( .Q(\SADR/m_fadrl[22] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgregadrh[22] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[20]  ( .Q(\SADR/m_fadrl[20] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgregadrh[20] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[17]  ( .Q(\SADR/m_fadrl[17] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[17] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[13]  ( .Q(\SADR/m_fadrl[13] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[13] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[18]  ( .Q(\SADR/m_fadrl[18] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgregadrh[18] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[11]  ( .Q(\SADR/m_fadrl[11] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[11] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[15]  ( .Q(\SADR/m_fadrl[15] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[15] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_invx1 \SADR/ADRFF/U150  ( .ZN(\SADR/ADRFF/n9120 ), .A(
        \SADR/ADRFF/n9119 ) );
    snl_invx1 \SADR/ADRFF/U152  ( .ZN(\SADR/ADRFF/n9122 ), .A(ad_latch) );
    snl_sffqenrnx1 \SADR/ADRFF/pgbitnoh_reg[0]  ( .Q(\pgbitnoh[0] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/intbitno[0] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgbitnoh_reg[1]  ( .Q(\pgbitnoh[1] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/intbitno[1] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[14]  ( .Q(\SADR/m_fadrl[14] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[14] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_invx1 \SADR/ADRFF/U151  ( .ZN(\SADR/ADRFF/n9121 ), .A(
        \SADR/ADRFF/n9119 ) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[26]  ( .Q(\pgsadrh[26] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[26] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[24]  ( .Q(\pgsadrh[24] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[24] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[17]  ( .Q(\pgsadrh[17] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[17] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[8]  ( .Q(\pgsadrh[8] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprlh[11] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgbitnoh_reg[3]  ( .Q(\pgbitnoh[3] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/intbitno[3] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[23]  ( .Q(\SADR/m_fadrl[23] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgregadrh[23] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[21]  ( .Q(\SADR/m_fadrl[21] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgregadrh[21] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[19]  ( .Q(\SADR/m_fadrl[19] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgregadrh[19] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[10]  ( .Q(\SADR/m_fadrl[10] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[10] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[12]  ( .Q(\SADR/m_fadrl[12] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[12] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrh_reg[31]  ( .Q(\SADR/m_fadrh[31] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprhh[31] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrh_reg[28]  ( .Q(\SADR/m_fadrh[28] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\pgsdprhh[28] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[16]  ( .Q(\SADR/m_fadrl[16] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[16] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[1]  ( .Q(\pgsadrh[1] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgsdprlh[4] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[5]  ( .Q(\SADR/m_fadrl[5] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[5] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[22]  ( .Q(\pgsadrh[22] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[22] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[20]  ( .Q(\pgsadrh[20] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[20] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[13]  ( .Q(\pgsadrh[13] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[13] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[11]  ( .Q(\pgsadrh[11] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[11] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[7]  ( .Q(\pgsadrh[7] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgsdprlh[10] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[5]  ( .Q(\pgsadrh[5] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgsdprlh[8] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[8]  ( .Q(\SADR/m_fadrl[8] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[8] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[18]  ( .Q(\pgsadrh[18] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9121 ), .SD(\SADR/sadr[18] ), .SE(
        \SADR/ADRFF/n9124 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[15]  ( .Q(\pgsadrh[15] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\SADR/sadr[15] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/pgsadrh_reg[3]  ( .Q(\pgsadrh[3] ), .D(1'b0), 
        .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgsdprlh[6] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_sffqenrnx1 \SADR/ADRFF/m_fadrl_reg[7]  ( .Q(\SADR/m_fadrl[7] ), .D(
        1'b0), .EN(1'b1), .RN(\SADR/ADRFF/n9120 ), .SD(\pgregadrh[7] ), .SE(
        \SADR/ADRFF/n9123 ), .CP(SCLK) );
    snl_and23x0 \REGF/pbmemff31/U166  ( .Z(\REGF/pbmemff31/RO_PSTA3B212[1] ), 
        .A(\pk_rwrit_h[56] ), .B(\pk_rwrit_h[48] ), .C(
        \REGF/pbmemff31/DO_SACONS ) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[19]  ( .Q(\REGF/RO_PCON[19] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[19]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[23]  ( .Q(\REGF/RO_PCON[23] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[23]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[10]  ( .Q(\REGF/RO_PCON[10] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[10]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[5]  ( .Q(\REGF/RO_PCON[5] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[5]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_invx05 \REGF/pbmemff31/U162  ( .ZN(\REGF/pbmemff31/n5647 ), .A(
        \REGF/n8052 ) );
    snl_invx05 \REGF/pbmemff31/U165  ( .ZN(\REGF/pbmemff31/n6437 ), .A(
        \pk_rwrit_h[56] ) );
    snl_and02x1 \REGF/pbmemff31/U167  ( .Z(\REGF/pbmemff31/RO_PSTA3B212[0] ), 
        .A(\REGF/pk_sctio_h ), .B(\REGF/pbmemff31/n5650 ) );
    snl_and02x1 \REGF/pbmemff31/U168  ( .Z(\REGF/pbmemff31/RO_EST13B291[2] ), 
        .A(ph_cperr_h), .B(\REGF/pbmemff31/n5651 ) );
    snl_nand12x1 \REGF/pbmemff31/U174  ( .ZN(\REGF/pbmemff31/n_729 ), .A(
        ph_stregwt_h), .B(\REGF/pbmemff31/n5651 ) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[8]  ( .Q(\REGF/RO_PCON[8] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[8]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[27]  ( .Q(\REGF/RO_PCON[27] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[27]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[1]  ( .Q(\REGF/RO_PCON[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[1]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PSTA3B_reg[1]  ( .Q(\REGF/RO_PSTA[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(
        \REGF/pbmemff31/RO_PSTA3B212[1] ), .SE(
        \REGF/pbmemff31/*cell*5410/U9/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[14]  ( .Q(\REGF/RO_PCON[14] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[14]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[3]  ( .Q(\REGF/RO_PCON[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[3]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_DTFLL_reg  ( .Q(\REGF/RO_EST2[15] ), .D(
        1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(\REGF/D2_DTFL ), 
        .SE(\REGF/pbmemff31/*cell*5410/U2/CONTROL1 ), .CP(SCLK) );
    snl_and02x1 \REGF/pbmemff31/U169  ( .Z(\REGF/pbmemff31/RO_EST13B291[1] ), 
        .A(ph_aluovf_h), .B(\REGF/pbmemff31/n5651 ) );
    snl_nor02x1 \REGF/pbmemff31/U172  ( .ZN(\REGF/pbmemff31/n5652 ), .A(
        ph_ex2regwt_h), .B(ph_stregwt_h) );
    snl_nand02x1 \REGF/pbmemff31/U173  ( .ZN(
        \REGF/pbmemff31/*cell*5410/U10/CONTROL1 ), .A(\REGF/pbmemff31/n5652 ), 
        .B(\REGF/pbmemff31/n5650 ) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[25]  ( .Q(\REGF/RO_PCON[25] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[25]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[16]  ( .Q(\REGF/RO_PCON[16] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[16]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[31]  ( .Q(pk_pcon31_h), .D(1'b0
        ), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[31]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[21]  ( .Q(\REGF/RO_PCON[21] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[21]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[12]  ( .Q(\REGF/RO_PCON[12] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[12]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[7]  ( .Q(\REGF/RO_PCON[7] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[7]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_EST13B_reg[1]  ( .Q(\REGF/RO_EST1[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(
        \REGF/pbmemff31/RO_EST13B291[1] ), .SE(\REGF/pbmemff31/n_729 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[28]  ( .Q(\REGF/RO_PCON[28] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[28]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_invx05 \REGF/pbmemff31/U175  ( .ZN(\REGF/pbmemff31/n5650 ), .A(
        \pk_rwrit_h[2] ) );
    snl_and02x1 \REGF/pbmemff31/U170  ( .Z(\REGF/pbmemff31/RO_EST13B291[0] ), 
        .A(pk_pcovf_h), .B(\REGF/pbmemff31/n5651 ) );
    snl_invx05 \REGF/pbmemff31/U177  ( .ZN(
        \REGF/pbmemff31/*cell*5410/U2/CONTROL1 ), .A(\REGF/pbmemff31/n5652 )
         );
    snl_or04x1 \REGF/pbmemff31/U171  ( .Z(
        \REGF/pbmemff31/*cell*5410/U9/CONTROL1 ), .A(ph_trsc_h), .B(
        \pk_rwrit_h[48] ), .C(\pk_rwrit_h[56] ), .D(ph_stregwt_h) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[20]  ( .Q(\REGF/RO_PCON[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[20]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[13]  ( .Q(\REGF/RO_PCON[13] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[13]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[6]  ( .Q(\REGF/RO_PCON[6] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[6]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_EST13B_reg[0]  ( .Q(\REGF/RO_EST1[1] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(
        \REGF/pbmemff31/RO_EST13B291[0] ), .SE(\REGF/pbmemff31/n_729 ), .CP(
        SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[30]  ( .Q(\REGF/RO_PCON[30] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[30]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[29]  ( .Q(\REGF/RO_PCON[29] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[29]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PEXE1B_reg  ( .Q(pk_pexe01_h), .D(1'b0), 
        .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[57] ), .CP(SCLK) );
    snl_invx1 \REGF/pbmemff31/U163  ( .ZN(\REGF/pbmemff31/n5648 ), .A(
        \REGF/pbmemff31/n5647 ) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[24]  ( .Q(\REGF/RO_PCON[24] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[24]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[2]  ( .Q(\REGF/RO_PCON[2] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[2]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[17]  ( .Q(\REGF/RO_PCON[17] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[17]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PSTA3B_reg[2]  ( .Q(\REGF/RO_PSTA[22] ), 
        .D(1'b0), .EN(\REGF/pbmemff31/n6437 ), .RN(\REGF/pbmemff31/n5648 ), 
        .SD(ph_pccons_h), .SE(ph_stregwt_h), .CP(SCLK) );
    snl_invx1 \REGF/pbmemff31/U164  ( .ZN(\REGF/pbmemff31/n5649 ), .A(
        \REGF/pbmemff31/n5647 ) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[9]  ( .Q(\REGF/RO_PCON[9] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[9]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PSTA3B_reg[0]  ( .Q(\REGF/RO_PSTA[20] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(
        \REGF/pbmemff31/RO_PSTA3B212[0] ), .SE(
        \REGF/pbmemff31/*cell*5410/U10/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \REGF/pbmemff31/U176  ( .ZN(\REGF/pbmemff31/n5651 ), .A(
        \pk_rwrit_h[55] ) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[26]  ( .Q(\REGF/RO_PCON[26] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[26]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[0]  ( .Q(\REGF/RO_PCON[0] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[0]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[18]  ( .Q(\REGF/RO_PCON[18] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[18]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[15]  ( .Q(\REGF/RO_PCON[15] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[15]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[22]  ( .Q(\REGF/RO_PCON[22] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(PDLIN[22]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[11]  ( .Q(\REGF/RO_PCON[11] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[11]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_PCON_reg[4]  ( .Q(\REGF/RO_PCON[4] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5649 ), .SD(PDLIN[4]), .SE(
        \pk_rwrit_h[58] ), .CP(SCLK) );
    snl_sffqenrnx1 \REGF/pbmemff31/RO_EST13B_reg[2]  ( .Q(\REGF/RO_EST1[3] ), 
        .D(1'b0), .EN(1'b1), .RN(\REGF/pbmemff31/n5648 ), .SD(
        \REGF/pbmemff31/RO_EST13B291[2] ), .SE(\REGF/pbmemff31/n_729 ), .CP(
        SCLK) );
    snl_ao012x1 \SAEXE/SRCRD/U29  ( .Z(\SAEXE/SRCRD/nrst[0] ), .A(
        \SAEXE/SRCRD/n93 ), .B(\SAEXE/SRCRD/erst[0] ), .C(\SAEXE/sa_start1 )
         );
    snl_ffqrnx1 \SAEXE/SRCRD/erst_reg[0]  ( .Q(\SAEXE/SRCRD/erst[0] ), .D(
        \SAEXE/SRCRD/nrst[0] ), .RN(n10735), .CP(SCLK) );
    snl_and02x1 \SAEXE/SRCRD/U30  ( .Z(\SAEXE/bnolth ), .A(
        \SAEXE/SRCRD/erst[0] ), .B(ph_lbend) );
    snl_invx05 \SAEXE/SRCRD/U32  ( .ZN(\SAEXE/SRCRD/n93 ), .A(ph_lbend) );
    snl_and23x0 \SAEXE/SRCRD/U31  ( .Z(\SAEXE/sa_start1 ), .A(
        \SAEXE/SRCRD/erst[0] ), .B(\SAEXE/exec_end1 ), .C(\SAEXE/srcrd_st ) );
    snl_ffqrnx1 \SAEXE/SRCRD/erst_reg[1]  ( .Q(\SAEXE/exec_end1 ), .D(
        \SAEXE/bnolth ), .RN(n10735), .CP(SCLK) );
    snl_muxi21x1 \ALUSHT/ALU/U364  ( .ZN(\ALUSHT/ALU/n2042 ), .A(
        \ALUSHT/ALU/n2140 ), .B(\ALUSHT/ALU/n2135 ), .S(\pgaluina[14] ) );
    snl_muxi21x1 \ALUSHT/ALU/U371  ( .ZN(\ALUSHT/ALU/n2026 ), .A(
        \ALUSHT/ALU/n2180 ), .B(\ALUSHT/ALU/n2181 ), .S(\pgaluina[2] ) );
    snl_aoi012x1 \ALUSHT/ALU/U394  ( .ZN(\ALUSHT/ALU/n1808 ), .A(
        \pgaluina[26] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U415  ( .ZN(\ALUSHT/ALU/n1830 ), .A(
        \pgaluinb[21] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U432  ( .ZN(\ALUSHT/ALU/pkaddina[20] ), .A(
        \ALUSHT/ALU/n1814 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nand02x1 \ALUSHT/ALU/U692  ( .ZN(\ALUSHT/ALU/n2242 ), .A(
        \ALUSHT/ALU/n2243 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nand02x1 \ALUSHT/ALU/U840  ( .ZN(\ALUSHT/ALU/n1819 ), .A(
        \ALUSHT/ALU/n2084 ), .B(\ALUSHT/ALU/n2083 ) );
    snl_muxi21x1 \ALUSHT/ALU/U702  ( .ZN(\ALUSHT/ALU/pkaddinb[8] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[8] ) );
    snl_muxi21x1 \ALUSHT/ALU/U725  ( .ZN(\ALUSHT/ALU/pkaddinb[16] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\ALUSHT/ALU/intb[16] )
         );
    snl_nand04x0 \ALUSHT/ALU/U529  ( .ZN(\ALUSHT/pkaluout[16] ), .A(
        \ALUSHT/ALU/n1970 ), .B(\ALUSHT/ALU/n1971 ), .C(\ALUSHT/ALU/n1972 ), 
        .D(\ALUSHT/ALU/n1973 ) );
    snl_invx05 \ALUSHT/ALU/U585  ( .ZN(\ALUSHT/ALU/n1852 ), .A(\pgaluina[1] )
         );
    snl_invx05 \ALUSHT/ALU/U867  ( .ZN(\ALUSHT/ALU/inta[29] ), .A(
        \ALUSHT/ALU/n1805 ) );
    snl_invx05 \ALUSHT/ALU/U560  ( .ZN(\ALUSHT/ALU/n1817 ), .A(\poalufnc[1] )
         );
    snl_xor3x1 \ALUSHT/ALU/U619  ( .Z(\ALUSHT/ALU/n2070 ), .A(
        \ALUSHT/ALU/n1906 ), .B(\ALUSHT/ALU/n2116 ), .C(\ALUSHT/ALU/n2117 ) );
    snl_xor2x0 \ALUSHT/ALU/U1047  ( .Z(\ALUSHT/ALU/n2112 ), .A(
        \ALUSHT/ALU/intb[21] ), .B(\ALUSHT/ALU/n1831 ) );
    snl_oai012x1 \ALUSHT/ALU/U650  ( .ZN(\ALUSHT/ALU/n2180 ), .A(\pgaluinb[2] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_ao022x1 \ALUSHT/ALU/U789  ( .Z(\ALUSHT/ALU/n2274 ), .A(
        \ALUSHT/ALU/pkdecout[23] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[23] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_nor02x2 \ALUSHT/ALU/U378  ( .ZN(\ALUSHT/ALU/n2095 ), .A(
        \ALUSHT/ALU/n2094 ), .B(\ALUSHT/ALU/n2075 ) );
    snl_nor02x1 \ALUSHT/ALU/U429  ( .ZN(\ALUSHT/ALU/pkaddina[23] ), .A(
        \ALUSHT/ALU/n1811 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U447  ( .ZN(\ALUSHT/ALU/pkaddina[4] ), .A(
        \ALUSHT/ALU/n1849 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor03x0 \ALUSHT/ALU/U547  ( .ZN(pkalucmf), .A(\ALUSHT/ALU/n2043 ), .B(
        \ALUSHT/ALU/n2044 ), .C(\ALUSHT/ALU/n2045 ) );
    snl_invx05 \ALUSHT/ALU/U882  ( .ZN(\ALUSHT/ALU/inta[25] ), .A(
        \ALUSHT/ALU/n1809 ) );
    snl_nor02x1 \ALUSHT/ALU/U912  ( .ZN(\ALUSHT/ALU/n1874 ), .A(
        \ALUSHT/ALU/n1835 ), .B(\ALUSHT/ALU/inta[16] ) );
    snl_nand02x1 \ALUSHT/ALU/U677  ( .ZN(\ALUSHT/ALU/n2220 ), .A(
        \ALUSHT/ALU/n2221 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U935  ( .ZN(\ALUSHT/ALU/n2004 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[8] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1029  ( .ZN(\ALUSHT/ALU/n1982 ), .A(
        \ALUSHT/ALU/n2238 ), .B(\ALUSHT/ALU/n2239 ), .S(\pgaluina[13] ) );
    snl_ao022x1 \ALUSHT/ALU/U777  ( .Z(\ALUSHT/ALU/n2268 ), .A(
        \ALUSHT/ALU/pkdecout[29] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[29] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_ao022x1 \ALUSHT/ALU/U809  ( .Z(\ALUSHT/ALU/n2283 ), .A(
        \ALUSHT/ALU/pkdecout[14] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[14] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U999  ( .ZN(\ALUSHT/ALU/n1952 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1830 ) );
    snl_oai222x0 \ALUSHT/ALU/U460  ( .ZN(\ALUSHT/ALU/pkincin[23] ), .A(
        \ALUSHT/ALU/n1828 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1811 ), .E(\ALUSHT/ALU/n1867 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_invx05 \ALUSHT/ALU/U835  ( .ZN(\ALUSHT/ALU/n2152 ), .A(
        \ALUSHT/ALU/n2055 ) );
    snl_nor02x1 \ALUSHT/ALU/U485  ( .ZN(\ALUSHT/ALU/pkdecin[29] ), .A(
        \ALUSHT/ALU/n1805 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nor04x0 \ALUSHT/ALU/U750  ( .ZN(\ALUSHT/ALU/n2050 ), .A(
        \ALUSHT/ALU/n1834 ), .B(\ALUSHT/ALU/n1835 ), .C(\ALUSHT/ALU/n2085 ), 
        .D(\ALUSHT/ALU/n2091 ) );
    snl_aoi112x0 \ALUSHT/ALU/U812  ( .ZN(\ALUSHT/ALU/n1985 ), .A(
        \ALUSHT/ALU/pkaddsum[13] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2284 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U982  ( .ZN(\ALUSHT/ALU/n1934 ), .A(
        \ALUSHT/ALU/n2195 ), .B(\ALUSHT/ALU/n2196 ), .S(\ALUSHT/ALU/inta[25] )
         );
    snl_nor02x1 \ALUSHT/ALU/U899  ( .ZN(\ALUSHT/ALU/n1870 ), .A(
        \ALUSHT/ALU/n1831 ), .B(\ALUSHT/ALU/inta[20] ) );
    snl_nor02x1 \ALUSHT/ALU/U909  ( .ZN(\ALUSHT/ALU/n1873 ), .A(
        \ALUSHT/ALU/n1834 ), .B(\ALUSHT/ALU/inta[17] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1015  ( .ZN(\ALUSHT/ALU/n2224 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[17] )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1032  ( .ZN(\ALUSHT/ALU/n1987 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1883 ) );
    snl_nand04x0 \ALUSHT/ALU/U515  ( .ZN(\ALUSHT/pkaluout[30] ), .A(
        \ALUSHT/ALU/n1914 ), .B(\ALUSHT/ALU/n1915 ), .C(\ALUSHT/ALU/n1916 ), 
        .D(\ALUSHT/ALU/n1917 ) );
    snl_nand04x0 \ALUSHT/ALU/U532  ( .ZN(\ALUSHT/pkaluout[13] ), .A(
        \ALUSHT/ALU/n1982 ), .B(\ALUSHT/ALU/n1983 ), .C(\ALUSHT/ALU/n1984 ), 
        .D(\ALUSHT/ALU/n1985 ) );
    snl_nand02x1 \ALUSHT/ALU/U602  ( .ZN(\ALUSHT/ALU/n2081 ), .A(
        \ALUSHT/ALU/n2090 ), .B(\ALUSHT/ALU/n2077 ) );
    snl_oa022x1 \ALUSHT/ALU/U625  ( .Z(\ALUSHT/ALU/n2123 ), .A(
        \ALUSHT/ALU/n2085 ), .B(\ALUSHT/ALU/n2124 ), .C(\ALUSHT/ALU/n2081 ), 
        .D(\pgaluina[15] ) );
    snl_muxi21x1 \ALUSHT/ALU/U967  ( .ZN(\ALUSHT/ALU/n1920 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1822 ) );
    snl_aoi112x0 \ALUSHT/ALU/U792  ( .ZN(\ALUSHT/ALU/n1949 ), .A(
        \ALUSHT/ALU/pkaddsum[22] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2275 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_oai012x1 \ALUSHT/ALU/U689  ( .ZN(\ALUSHT/ALU/n2238 ), .A(
        \pgaluinb[13] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U940  ( .ZN(\ALUSHT/ALU/n2011 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1895 ) );
    snl_muxi21x1 \ALUSHT/ALU/U719  ( .ZN(\ALUSHT/ALU/pkaddinb[21] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1830 ) );
    snl_nor02x1 \ALUSHT/ALU/U497  ( .ZN(\ALUSHT/ALU/pkdecin[17] ), .A(
        \ALUSHT/ALU/n1837 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_and02x1 \ALUSHT/ALU/U507  ( .Z(\ALUSHT/ALU/pkdecin[6] ), .A(
        \pgaluina[6] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_invx05 \ALUSHT/ALU/U849  ( .ZN(\ALUSHT/ALU/n2090 ), .A(
        \ALUSHT/ALU/n2048 ) );
    snl_muxi21x1 \ALUSHT/ALU/U975  ( .ZN(\ALUSHT/ALU/n1928 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1824 ) );
    snl_nand04x0 \ALUSHT/ALU/U520  ( .ZN(\ALUSHT/pkaluout[25] ), .A(
        \ALUSHT/ALU/n1934 ), .B(\ALUSHT/ALU/n1935 ), .C(\ALUSHT/ALU/n1936 ), 
        .D(\ALUSHT/ALU/n1937 ) );
    snl_nand02x1 \ALUSHT/ALU/U610  ( .ZN(\ALUSHT/ALU/n2046 ), .A(
        \ALUSHT/ALU/n2092 ), .B(\ALUSHT/ALU/n2073 ) );
    snl_oai012x1 \ALUSHT/ALU/U637  ( .ZN(\ALUSHT/ALU/n2160 ), .A(\pgaluinb[6] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_aoi112x0 \ALUSHT/ALU/U780  ( .ZN(\ALUSHT/ALU/n1925 ), .A(
        \ALUSHT/ALU/pkaddsum[28] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2269 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U952  ( .ZN(\ALUSHT/ALU/n2024 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[3] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1007  ( .ZN(\ALUSHT/ALU/n2218 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1832 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1020  ( .ZN(\ALUSHT/ALU/n1971 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1874 ) );
    snl_oai012x2 \ALUSHT/ALU/U381  ( .ZN(\ALUSHT/ALU/n2143 ), .A(
        \ALUSHT/ALU/n2079 ), .B(\ALUSHT/ALU/n2046 ), .C(\ALUSHT/ALU/n2144 ) );
    snl_ao022x4 \ALUSHT/ALU/U386  ( .Z(\ALUSHT/ALU/n2267 ), .A(
        \ALUSHT/ALU/pkdecout[2] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[2] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_aoi012x1 \ALUSHT/ALU/U407  ( .ZN(\ALUSHT/ALU/n1822 ), .A(
        \pgaluinb[29] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_aoi012x1 \ALUSHT/ALU/U420  ( .ZN(\ALUSHT/ALU/n1835 ), .A(
        \pgaluinb[16] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_oai222x0 \ALUSHT/ALU/U455  ( .ZN(\ALUSHT/ALU/pkincin[28] ), .A(
        \ALUSHT/ALU/n1823 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1806 ), .E(\ALUSHT/ALU/n1862 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_invx05 \ALUSHT/ALU/U569  ( .ZN(\ALUSHT/ALU/n1890 ), .A(\pgaluinb[8] )
         );
    snl_nand02x1 \ALUSHT/ALU/U659  ( .ZN(\ALUSHT/ALU/n2193 ), .A(
        \ALUSHT/ALU/n2194 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_aoi112x0 \ALUSHT/ALU/U765  ( .ZN(\ALUSHT/ALU/n2013 ), .A(
        \ALUSHT/ALU/pkaddsum[6] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2261 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_xnor2x0 \ALUSHT/ALU/U827  ( .ZN(\ALUSHT/ALU/n2071 ), .A(
        \ALUSHT/ALU/n1902 ), .B(\pgaluinb[1] ) );
    snl_oai222x0 \ALUSHT/ALU/U469  ( .ZN(\ALUSHT/ALU/pkincin[14] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1878 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1839 ), .E(\ALUSHT/ALU/n1879 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai222x0 \ALUSHT/ALU/U472  ( .ZN(\ALUSHT/ALU/pkincin[11] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1884 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1842 ), .E(\ALUSHT/ALU/n1885 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_aoi112x0 \ALUSHT/ALU/U800  ( .ZN(\ALUSHT/ALU/n1961 ), .A(
        \ALUSHT/ALU/pkaddsum[19] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2279 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U990  ( .ZN(\ALUSHT/ALU/n1942 ), .A(
        \ALUSHT/ALU/n2201 ), .B(\ALUSHT/ALU/n2202 ), .S(\ALUSHT/ALU/inta[23] )
         );
    snl_nor04x0 \ALUSHT/ALU/U742  ( .ZN(\ALUSHT/ALU/n2089 ), .A(
        \ALUSHT/ALU/n1888 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1890 ), 
        .D(\ALUSHT/ALU/n1892 ) );
    snl_aoi112x0 \ALUSHT/ALU/U759  ( .ZN(\ALUSHT/ALU/n2001 ), .A(
        \ALUSHT/ALU/pkaddsum[9] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2258 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_xor3x1 \ALUSHT/ALU/U555  ( .Z(\ALUSHT/ALU/n2047 ), .A(
        \ALUSHT/ALU/n2070 ), .B(\ALUSHT/ALU/n2071 ), .C(\ALUSHT/ALU/n2072 ) );
    snl_invx05 \ALUSHT/ALU/U572  ( .ZN(\ALUSHT/ALU/n1847 ), .A(\pgaluina[6] )
         );
    snl_nand02x1 \ALUSHT/ALU/U642  ( .ZN(\ALUSHT/ALU/n2167 ), .A(
        \ALUSHT/ALU/n2168 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nor02x1 \ALUSHT/ALU/U890  ( .ZN(\ALUSHT/ALU/n1867 ), .A(
        \ALUSHT/ALU/n1828 ), .B(\ALUSHT/ALU/inta[23] ) );
    snl_nor02x1 \ALUSHT/ALU/U900  ( .ZN(\ALUSHT/ALU/n1905 ), .A(
        \ALUSHT/ALU/n1904 ), .B(\pgaluina[1] ) );
    snl_muxi21x1 \ALUSHT/ALU/U927  ( .ZN(\ALUSHT/ALU/n2141 ), .A(
        \ALUSHT/ALU/n2134 ), .B(\ALUSHT/ALU/n2130 ), .S(\ALUSHT/ALU/n1803 ) );
    snl_nand02x1 \ALUSHT/ALU/U665  ( .ZN(\ALUSHT/ALU/n2202 ), .A(
        \ALUSHT/ALU/n2203 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nor02x1 \ALUSHT/ALU/U852  ( .ZN(\ALUSHT/ALU/n1891 ), .A(
        \ALUSHT/ALU/n1890 ), .B(\pgaluina[8] ) );
    snl_muxi21x1 \ALUSHT/ALU/U949  ( .ZN(\ALUSHT/ALU/n2020 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[4] ) );
    snl_invx05 \ALUSHT/ALU/U597  ( .ZN(\ALUSHT/ALU/n1853 ), .A(\pgaluina[0] )
         );
    snl_oai012x1 \ALUSHT/ALU/U680  ( .ZN(\ALUSHT/ALU/n2225 ), .A(
        \ALUSHT/ALU/intb[16] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U710  ( .ZN(\ALUSHT/ALU/pkaddinb[2] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1902 ) );
    snl_or08x1 \ALUSHT/ALU/U737  ( .Z(\ALUSHT/ALU/n2038 ), .A(
        \ALUSHT/ALU/n1860 ), .B(\ALUSHT/ALU/n2118 ), .C(\ALUSHT/ALU/n1887 ), 
        .D(\ALUSHT/ALU/n1907 ), .E(\ALUSHT/ALU/n1883 ), .F(\ALUSHT/ALU/n1885 ), 
        .G(\ALUSHT/ALU/n1879 ), .H(\ALUSHT/ALU/n1881 ) );
    snl_invx05 \ALUSHT/ALU/U875  ( .ZN(\ALUSHT/ALU/inta[27] ), .A(
        \ALUSHT/ALU/n1807 ) );
    snl_muxi21x1 \ALUSHT/ALU/U969  ( .ZN(\ALUSHT/ALU/n1923 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1862 ) );
    snl_xnor2x0 \ALUSHT/ALU/U1052  ( .ZN(\ALUSHT/ALU/n2116 ), .A(
        \ALUSHT/ALU/n1890 ), .B(\ALUSHT/ALU/n1886 ) );
    snl_aoi012x1 \ALUSHT/ALU/U400  ( .ZN(\ALUSHT/ALU/n1814 ), .A(
        \pgaluina[20] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nor02x1 \ALUSHT/ALU/U427  ( .ZN(\ALUSHT/ALU/pkaddina[25] ), .A(
        \ALUSHT/ALU/n1809 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_invx05 \ALUSHT/ALU/U590  ( .ZN(\ALUSHT/ALU/n1880 ), .A(\pgaluinb[13] )
         );
    snl_oai012x1 \ALUSHT/ALU/U687  ( .ZN(\ALUSHT/ALU/n2235 ), .A(
        \pgaluinb[14] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U730  ( .ZN(\ALUSHT/ALU/pkaddinb[10] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[10] ) );
    snl_invx05 \ALUSHT/ALU/U872  ( .ZN(\ALUSHT/ALU/intb[28] ), .A(
        \ALUSHT/ALU/n1823 ) );
    snl_muxi21x1 \ALUSHT/ALU/U717  ( .ZN(\ALUSHT/ALU/pkaddinb[23] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1828 ) );
    snl_nor02x1 \ALUSHT/ALU/U449  ( .ZN(\ALUSHT/ALU/pkaddina[2] ), .A(
        \ALUSHT/ALU/n1851 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_ao022x1 \ALUSHT/ALU/U779  ( .Z(\ALUSHT/ALU/n2269 ), .A(
        \ALUSHT/ALU/pkdecout[28] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[28] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_nor02x1 \ALUSHT/ALU/U855  ( .ZN(\ALUSHT/ALU/n1897 ), .A(
        \ALUSHT/ALU/n1896 ), .B(\pgaluina[5] ) );
    snl_and08x1 \ALUSHT/ALU/U552  ( .Z(\ALUSHT/ALU/n2058 ), .A(
        \ALUSHT/ALU/n2059 ), .B(\ALUSHT/ALU/n2060 ), .C(\ALUSHT/ALU/n2061 ), 
        .D(\ALUSHT/ALU/n2062 ), .E(\ALUSHT/ALU/n2063 ), .F(\ALUSHT/ALU/n2064 ), 
        .G(\ALUSHT/ALU/n2065 ), .H(\ALUSHT/ALU/n2066 ) );
    snl_oai012x1 \ALUSHT/ALU/U662  ( .ZN(\ALUSHT/ALU/n2198 ), .A(
        \ALUSHT/ALU/intb[24] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_invx05 \ALUSHT/ALU/U575  ( .ZN(\ALUSHT/ALU/n1896 ), .A(\pgaluinb[5] )
         );
    snl_invx05 \ALUSHT/ALU/U920  ( .ZN(\ALUSHT/ALU/n2230 ), .A(
        \ALUSHT/ALU/n2153 ) );
    snl_muxi21x1 \ALUSHT/ALU/U365  ( .ZN(\ALUSHT/ALU/n2034 ), .A(
        \ALUSHT/ALU/n2250 ), .B(\ALUSHT/ALU/n2251 ), .S(\pgaluina[0] ) );
    snl_nand02x2 \ALUSHT/ALU/U376  ( .ZN(\ALUSHT/ALU/n2151 ), .A(
        \ALUSHT/ALU/n2099 ), .B(\ALUSHT/ALU/n2152 ) );
    snl_aoi0b12x2 \ALUSHT/ALU/U388  ( .ZN(\ALUSHT/ALU/n2148 ), .A(
        \ALUSHT/ALU/n2083 ), .B(\ALUSHT/ALU/n2096 ), .C(\ALUSHT/ALU/n2144 ) );
    snl_ao0b12x1 \ALUSHT/ALU/U452  ( .Z(\ALUSHT/ALU/pkincin[31] ), .A(
        \ALUSHT/ALU/n1854 ), .B(\ALUSHT/ALU/n1855 ), .C(\ALUSHT/ALU/n1856 ) );
    snl_oai222x0 \ALUSHT/ALU/U475  ( .ZN(\ALUSHT/ALU/pkincin[8] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1890 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1845 ), .E(\ALUSHT/ALU/n1891 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_aoi033x0 \ALUSHT/ALU/U549  ( .ZN(\ALUSHT/ALU/n2049 ), .A(
        \ALUSHT/ALU/n2050 ), .B(\ALUSHT/ALU/n2051 ), .C(\ALUSHT/ALU/n2052 ), 
        .D(\ALUSHT/ALU/pkcmpina[31] ), .E(\pgaluina[15] ), .F(
        \ALUSHT/ALU/n2053 ) );
    snl_oai012x1 \ALUSHT/ALU/U645  ( .ZN(\ALUSHT/ALU/n2172 ), .A(
        \ALUSHT/ALU/pkcmpinb[31] ), .B(\ALUSHT/ALU/n2146 ), .C(
        \ALUSHT/ALU/n2098 ) );
    snl_invx05 \ALUSHT/ALU/U897  ( .ZN(\ALUSHT/ALU/inta[20] ), .A(
        \ALUSHT/ALU/n1814 ) );
    snl_invx05 \ALUSHT/ALU/U907  ( .ZN(\ALUSHT/ALU/n1837 ), .A(
        \ALUSHT/ALU/inta[17] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1000  ( .ZN(\ALUSHT/ALU/n2212 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[20] )
         );
    snl_nand02x1 \ALUSHT/ALU/U679  ( .ZN(\ALUSHT/ALU/n2223 ), .A(
        \ALUSHT/ALU/n2224 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1027  ( .ZN(\ALUSHT/ALU/n2240 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[13] ) );
    snl_nor04x0 \ALUSHT/ALU/U745  ( .ZN(\ALUSHT/ALU/n2086 ), .A(
        \ALUSHT/ALU/n1882 ), .B(\ALUSHT/ALU/n1884 ), .C(\ALUSHT/ALU/n1886 ), 
        .D(\ALUSHT/ALU/n1906 ) );
    snl_aoi022x1 \ALUSHT/ALU/U807  ( .ZN(\ALUSHT/ALU/n1976 ), .A(
        \ALUSHT/ALU/pkincout[15] ), .B(\ALUSHT/ALU/n1855 ), .C(
        \ALUSHT/ALU/pkdecout[15] ), .D(\ALUSHT/ALU/n1909 ) );
    snl_muxi21x1 \ALUSHT/ALU/U997  ( .ZN(\ALUSHT/ALU/n1951 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1869 ) );
    snl_oai222x0 \ALUSHT/ALU/U482  ( .ZN(\ALUSHT/ALU/pkincin[1] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1904 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1852 ), .E(\ALUSHT/ALU/n1905 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nor02x1 \ALUSHT/ALU/U490  ( .ZN(\ALUSHT/ALU/pkdecin[24] ), .A(
        \ALUSHT/ALU/n1810 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand04x0 \ALUSHT/ALU/U527  ( .ZN(\ALUSHT/pkaluout[18] ), .A(
        \ALUSHT/ALU/n1962 ), .B(\ALUSHT/ALU/n1963 ), .C(\ALUSHT/ALU/n1964 ), 
        .D(\ALUSHT/ALU/n1965 ) );
    snl_ao022x1 \ALUSHT/ALU/U762  ( .Z(\ALUSHT/ALU/n2260 ), .A(
        \ALUSHT/ALU/pkdecout[7] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[7] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_aoi112x0 \ALUSHT/ALU/U820  ( .ZN(\ALUSHT/ALU/n2037 ), .A(
        \ALUSHT/ALU/pkaddsum[0] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2288 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U869  ( .ZN(\ALUSHT/ALU/n1861 ), .A(
        \ALUSHT/ALU/n1822 ), .B(\ALUSHT/ALU/inta[29] ) );
    snl_xor3x1 \ALUSHT/ALU/U617  ( .Z(\ALUSHT/ALU/n2109 ), .A(
        \ALUSHT/ALU/n2110 ), .B(\ALUSHT/ALU/n2111 ), .C(\ALUSHT/ALU/n2112 ) );
    snl_muxi21x1 \ALUSHT/ALU/U955  ( .ZN(\ALUSHT/ALU/n1910 ), .A(
        \ALUSHT/ALU/n2172 ), .B(\ALUSHT/ALU/n2173 ), .S(\ALUSHT/ALU/n1854 ) );
    snl_xnor2x0 \ALUSHT/ALU/U1049  ( .ZN(\ALUSHT/ALU/n2115 ), .A(
        \ALUSHT/ALU/n1875 ), .B(\ALUSHT/ALU/n1878 ) );
    snl_and08x1 \ALUSHT/ALU/U630  ( .Z(\ALUSHT/ALU/n2140 ), .A(
        \ALUSHT/ALU/n1851 ), .B(\ALUSHT/ALU/n1850 ), .C(\ALUSHT/ALU/n1849 ), 
        .D(\ALUSHT/ALU/n1848 ), .E(\ALUSHT/ALU/n1853 ), .F(\ALUSHT/ALU/n1852 ), 
        .G(\ALUSHT/ALU/n2141 ), .H(\ALUSHT/ALU/n2142 ) );
    snl_ao022x1 \ALUSHT/ALU/U787  ( .Z(\ALUSHT/ALU/n2273 ), .A(
        \ALUSHT/ALU/pkdecout[24] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[24] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_and02x1 \ALUSHT/ALU/U500  ( .Z(\ALUSHT/ALU/pkdecin[13] ), .A(
        \pgaluina[13] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_and02x1 \ALUSHT/ALU/U512  ( .Z(\ALUSHT/ALU/pkdecin[1] ), .A(
        \pgaluina[1] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_nand04x0 \ALUSHT/ALU/U535  ( .ZN(\ALUSHT/pkaluout[10] ), .A(
        \ALUSHT/ALU/n1994 ), .B(\ALUSHT/ALU/n1995 ), .C(\ALUSHT/ALU/n1996 ), 
        .D(\ALUSHT/ALU/n1997 ) );
    snl_muxi21x1 \ALUSHT/ALU/U947  ( .ZN(\ALUSHT/ALU/n2019 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1899 ) );
    snl_muxi21x1 \ALUSHT/ALU/U972  ( .ZN(\ALUSHT/ALU/n2191 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[27] )
         );
    snl_invx05 \ALUSHT/ALU/U605  ( .ZN(\ALUSHT/ALU/n2045 ), .A(\poalufnc[3] )
         );
    snl_ao022x1 \ALUSHT/ALU/U795  ( .Z(\ALUSHT/ALU/n2277 ), .A(
        \ALUSHT/ALU/pkdecout[20] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[20] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_nand12x1 \ALUSHT/ALU/U622  ( .ZN(\ALUSHT/ALU/n2120 ), .A(
        \ALUSHT/ALU/pkaddinb[15] ), .B(\ALUSHT/ALU/pkaddsum[15] ) );
    snl_muxi21x1 \ALUSHT/ALU/U960  ( .ZN(\ALUSHT/ALU/n1916 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1820 ) );
    snl_nand02x1 \ALUSHT/ALU/U599  ( .ZN(\ALUSHT/ALU/n2082 ), .A(\poalufnc[0] 
        ), .B(\ALUSHT/ALU/n1817 ) );
    snl_or04x1 \ALUSHT/ALU/U739  ( .Z(\ALUSHT/ALU/n2132 ), .A(
        \ALUSHT/ALU/inta[18] ), .B(\ALUSHT/ALU/inta[19] ), .C(
        \ALUSHT/ALU/inta[20] ), .D(\ALUSHT/ALU/inta[21] ) );
    snl_aoi012x1 \ALUSHT/ALU/U409  ( .ZN(\ALUSHT/ALU/n1824 ), .A(
        \pgaluinb[27] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U440  ( .ZN(\ALUSHT/ALU/pkaddina[11] ), .A(
        \ALUSHT/ALU/n1842 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U467  ( .ZN(\ALUSHT/ALU/pkincin[16] ), .A(
        \ALUSHT/ALU/n1835 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1838 ), .E(\ALUSHT/ALU/n1874 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nor04x0 \ALUSHT/ALU/U757  ( .ZN(\ALUSHT/ALU/n2136 ), .A(
        \ALUSHT/ALU/n1851 ), .B(\ALUSHT/ALU/n1852 ), .C(\ALUSHT/ALU/n1840 ), 
        .D(\ALUSHT/ALU/n1841 ) );
    snl_ao022x1 \ALUSHT/ALU/U815  ( .Z(\ALUSHT/ALU/n2286 ), .A(
        \ALUSHT/ALU/pkdecout[11] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[11] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U985  ( .ZN(\ALUSHT/ALU/n1939 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1866 ) );
    snl_nor02x1 \ALUSHT/ALU/U832  ( .ZN(\ALUSHT/ALU/n2233 ), .A(
        \ALUSHT/ALU/n2094 ), .B(\ALUSHT/ALU/n2048 ) );
    snl_nand04x0 \ALUSHT/ALU/U540  ( .ZN(\ALUSHT/pkaluout[5] ), .A(
        \ALUSHT/ALU/n2014 ), .B(\ALUSHT/ALU/n2015 ), .C(\ALUSHT/ALU/n2016 ), 
        .D(\ALUSHT/ALU/n2017 ) );
    snl_oai012x1 \ALUSHT/ALU/U670  ( .ZN(\ALUSHT/ALU/n2210 ), .A(
        \ALUSHT/ALU/intb[20] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_ao022x1 \ALUSHT/ALU/U770  ( .Z(\ALUSHT/ALU/n2264 ), .A(
        \ALUSHT/ALU/pkdecout[3] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[3] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U929  ( .ZN(\ALUSHT/ALU/n1999 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1889 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1012  ( .ZN(\ALUSHT/ALU/n1963 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1872 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1035  ( .ZN(\ALUSHT/ALU/n2246 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[11] ) );
    snl_muxi21x1 \ALUSHT/ALU/U932  ( .ZN(\ALUSHT/ALU/n2156 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1890 ) );
    snl_invx05 \ALUSHT/ALU/U885  ( .ZN(\ALUSHT/ALU/inta[24] ), .A(
        \ALUSHT/ALU/n1810 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1009  ( .ZN(\ALUSHT/ALU/n1958 ), .A(
        \ALUSHT/ALU/n2216 ), .B(\ALUSHT/ALU/n2217 ), .S(\ALUSHT/ALU/inta[19] )
         );
    snl_nor02x1 \ALUSHT/ALU/U915  ( .ZN(\ALUSHT/ALU/n1881 ), .A(
        \ALUSHT/ALU/n1880 ), .B(\pgaluina[13] ) );
    snl_aoi012x1 \ALUSHT/ALU/U393  ( .ZN(\ALUSHT/ALU/n1807 ), .A(
        \pgaluina[27] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nand02x1 \ALUSHT/ALU/U567  ( .ZN(\ALUSHT/ALU/n2079 ), .A(\poalufnc[0] 
        ), .B(\poalufnc[1] ) );
    snl_invx05 \ALUSHT/ALU/U582  ( .ZN(\ALUSHT/ALU/n1875 ), .A(\pgaluinb[15] )
         );
    snl_nand02x1 \ALUSHT/ALU/U657  ( .ZN(\ALUSHT/ALU/n2190 ), .A(
        \ALUSHT/ALU/n2191 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_invx05 \ALUSHT/ALU/U829  ( .ZN(\ALUSHT/ALU/n2124 ), .A(
        \ALUSHT/ALU/n2091 ) );
    snl_invx05 \ALUSHT/ALU/U860  ( .ZN(\ALUSHT/ALU/n2060 ), .A(
        \ALUSHT/ALU/pkcmpinb[31] ) );
    snl_aoi012x1 \ALUSHT/ALU/U412  ( .ZN(\ALUSHT/ALU/n1827 ), .A(
        \pgaluinb[24] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U435  ( .ZN(\ALUSHT/ALU/pkaddina[17] ), .A(
        \ALUSHT/ALU/n1837 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai012x1 \ALUSHT/ALU/U695  ( .ZN(\ALUSHT/ALU/n2247 ), .A(
        \pgaluinb[10] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U705  ( .ZN(\ALUSHT/ALU/pkaddinb[5] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[5] ) );
    snl_muxi21x1 \ALUSHT/ALU/U722  ( .ZN(\ALUSHT/ALU/pkaddinb[19] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1832 ) );
    snl_invx05 \ALUSHT/ALU/U847  ( .ZN(\ALUSHT/ALU/n2083 ), .A(
        \ALUSHT/ALU/n2082 ) );
    snl_nor02x1 \ALUSHT/ALU/U448  ( .ZN(\ALUSHT/ALU/pkaddina[3] ), .A(
        \ALUSHT/ALU/n1850 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U453  ( .ZN(\ALUSHT/ALU/pkincin[30] ), .A(
        \ALUSHT/ALU/n1820 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1802 ), .E(\ALUSHT/ALU/n1859 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai222x0 \ALUSHT/ALU/U474  ( .ZN(\ALUSHT/ALU/pkincin[9] ), .A(
        \ALUSHT/ALU/n1888 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1844 ), .E(\ALUSHT/ALU/n1889 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nor02x1 \ALUSHT/ALU/U491  ( .ZN(\ALUSHT/ALU/pkdecin[23] ), .A(
        \ALUSHT/ALU/n1811 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nor02x1 \ALUSHT/ALU/U499  ( .ZN(\ALUSHT/ALU/pkdecin[14] ), .A(
        \ALUSHT/ALU/n1839 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_and02x1 \ALUSHT/ALU/U509  ( .Z(\ALUSHT/ALU/pkdecin[4] ), .A(
        \pgaluina[4] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_and02x1 \ALUSHT/ALU/U501  ( .Z(\ALUSHT/ALU/pkdecin[12] ), .A(
        \pgaluina[12] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_nand04x0 \ALUSHT/ALU/U526  ( .ZN(\ALUSHT/pkaluout[19] ), .A(
        \ALUSHT/ALU/n1958 ), .B(\ALUSHT/ALU/n1959 ), .C(\ALUSHT/ALU/n1960 ), 
        .D(\ALUSHT/ALU/n1961 ) );
    snl_oai012x1 \ALUSHT/ALU/U639  ( .ZN(\ALUSHT/ALU/n2163 ), .A(\pgaluinb[5] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_invx05 \ALUSHT/ALU/U868  ( .ZN(\ALUSHT/ALU/intb[29] ), .A(
        \ALUSHT/ALU/n1822 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1040  ( .ZN(\ALUSHT/ALU/n1996 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[10] ) );
    snl_xor2x0 \ALUSHT/ALU/U1048  ( .Z(\ALUSHT/ALU/n2292 ), .A(
        \ALUSHT/ALU/intb[19] ), .B(\ALUSHT/ALU/n1833 ) );
    snl_xor3x1 \ALUSHT/ALU/U616  ( .Z(\ALUSHT/ALU/n2106 ), .A(
        \ALUSHT/ALU/intb[17] ), .B(\ALUSHT/ALU/n2107 ), .C(\ALUSHT/ALU/n2108 )
         );
    snl_aoi112x0 \ALUSHT/ALU/U786  ( .ZN(\ALUSHT/ALU/n1937 ), .A(
        \ALUSHT/ALU/pkaddsum[25] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2272 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U954  ( .ZN(\ALUSHT/ALU/n1911 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2233 ), .S(\ALUSHT/ALU/n2256 ) );
    snl_oai012x1 \ALUSHT/ALU/U631  ( .ZN(\ALUSHT/ALU/n2147 ), .A(\pgaluinb[9] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_nor03x0 \ALUSHT/ALU/U548  ( .ZN(pkaluopc), .A(\ALUSHT/ALU/n2046 ), .B(
        \ALUSHT/ALU/n2047 ), .C(\ALUSHT/ALU/n2048 ) );
    snl_muxi21x1 \ALUSHT/ALU/U973  ( .ZN(\ALUSHT/ALU/n1927 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1863 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1001  ( .ZN(\ALUSHT/ALU/n1955 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1870 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1026  ( .ZN(\ALUSHT/ALU/n1980 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[14] ) );
    snl_oai012x1 \ALUSHT/ALU/U678  ( .ZN(\ALUSHT/ALU/n2222 ), .A(
        \ALUSHT/ALU/intb[17] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_nor04x0 \ALUSHT/ALU/U744  ( .ZN(\ALUSHT/ALU/n2087 ), .A(
        \ALUSHT/ALU/n1902 ), .B(\ALUSHT/ALU/n1904 ), .C(\ALUSHT/ALU/n1878 ), 
        .D(\ALUSHT/ALU/n1880 ) );
    snl_aoi112x0 \ALUSHT/ALU/U806  ( .ZN(\ALUSHT/ALU/n1973 ), .A(
        \ALUSHT/ALU/pkaddsum[16] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2282 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U996  ( .ZN(\ALUSHT/ALU/n2209 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1830 ) );
    snl_aoi112x0 \ALUSHT/ALU/U763  ( .ZN(\ALUSHT/ALU/n2009 ), .A(
        \ALUSHT/ALU/pkaddsum[7] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2260 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_xor2x0 \ALUSHT/ALU/U821  ( .Z(\ALUSHT/ALU/n2289 ), .A(
        \ALUSHT/ALU/intb[27] ), .B(\ALUSHT/ALU/intb[26] ) );
    snl_aoi112x0 \ALUSHT/ALU/U778  ( .ZN(\ALUSHT/ALU/n1921 ), .A(
        \ALUSHT/ALU/pkaddsum[29] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2268 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U553  ( .ZN(\ALUSHT/ALU/n2067 ), .A(\poalufnc[1] ), 
        .B(\ALUSHT/ALU/n2068 ) );
    snl_nand02x1 \ALUSHT/ALU/U663  ( .ZN(\ALUSHT/ALU/n2199 ), .A(
        \ALUSHT/ALU/n2200 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_invx05 \ALUSHT/ALU/U921  ( .ZN(\ALUSHT/ALU/n2228 ), .A(
        \ALUSHT/ALU/n2145 ) );
    snl_oai012x2 \ALUSHT/ALU/U380  ( .ZN(\ALUSHT/ALU/n2153 ), .A(
        \ALUSHT/ALU/n2075 ), .B(\ALUSHT/ALU/n2046 ), .C(\ALUSHT/ALU/n2101 ) );
    snl_aoi012x1 \ALUSHT/ALU/U401  ( .ZN(\ALUSHT/ALU/n1815 ), .A(
        \pgaluina[19] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_invx05 \ALUSHT/ALU/U574  ( .ZN(\ALUSHT/ALU/n1848 ), .A(\pgaluina[5] )
         );
    snl_invx05 \ALUSHT/ALU/U591  ( .ZN(\ALUSHT/ALU/n1841 ), .A(\pgaluina[12] )
         );
    snl_nand02x1 \ALUSHT/ALU/U644  ( .ZN(\ALUSHT/ALU/n2170 ), .A(
        \ALUSHT/ALU/n2171 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nor02x1 \ALUSHT/ALU/U896  ( .ZN(\ALUSHT/ALU/n1869 ), .A(
        \ALUSHT/ALU/n1830 ), .B(\ALUSHT/ALU/inta[21] ) );
    snl_nor02x1 \ALUSHT/ALU/U906  ( .ZN(\ALUSHT/ALU/n1872 ), .A(
        \ALUSHT/ALU/n1833 ), .B(\ALUSHT/ALU/inta[18] ) );
    snl_muxi21x1 \ALUSHT/ALU/U968  ( .ZN(\ALUSHT/ALU/n2188 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[28] )
         );
    snl_xnor2x0 \ALUSHT/ALU/U1053  ( .ZN(\ALUSHT/ALU/n2117 ), .A(
        \ALUSHT/ALU/n1894 ), .B(\ALUSHT/ALU/n1892 ) );
    snl_aoi012x1 \ALUSHT/ALU/U392  ( .ZN(\ALUSHT/ALU/n1806 ), .A(
        \pgaluina[28] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U413  ( .ZN(\ALUSHT/ALU/n1828 ), .A(
        \pgaluinb[23] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U426  ( .ZN(\ALUSHT/ALU/pkaddina[26] ), .A(
        \ALUSHT/ALU/n1808 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_muxi21x1 \ALUSHT/ALU/U686  ( .ZN(\ALUSHT/ALU/n2234 ), .A(
        \ALUSHT/ALU/n2174 ), .B(\ALUSHT/ALU/n2146 ), .S(\ALUSHT/ALU/n1877 ) );
    snl_muxi21x1 \ALUSHT/ALU/U716  ( .ZN(\ALUSHT/ALU/pkaddinb[24] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1827 ) );
    snl_muxi21x1 \ALUSHT/ALU/U731  ( .ZN(\ALUSHT/ALU/pkaddinb[0] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[0] ) );
    snl_nor02x1 \ALUSHT/ALU/U873  ( .ZN(\ALUSHT/ALU/n1862 ), .A(
        \ALUSHT/ALU/inta[28] ), .B(\ALUSHT/ALU/n1823 ) );
    snl_nor02x1 \ALUSHT/ALU/U854  ( .ZN(\ALUSHT/ALU/n1895 ), .A(
        \ALUSHT/ALU/n1894 ), .B(\pgaluina[6] ) );
    snl_nand02x1 \ALUSHT/ALU/U861  ( .ZN(\ALUSHT/ALU/n1855 ), .A(
        \ALUSHT/ALU/n1858 ), .B(\ALUSHT/ALU/n1860 ) );
    snl_nor02x1 \ALUSHT/ALU/U434  ( .ZN(\ALUSHT/ALU/pkaddina[18] ), .A(
        \ALUSHT/ALU/n1816 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_invx05 \ALUSHT/ALU/U583  ( .ZN(\ALUSHT/ALU/n1851 ), .A(\pgaluina[2] )
         );
    snl_nand02x1 \ALUSHT/ALU/U694  ( .ZN(\ALUSHT/ALU/n2245 ), .A(
        \ALUSHT/ALU/n2246 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U723  ( .ZN(\ALUSHT/ALU/pkaddinb[18] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1833 ) );
    snl_muxi21x1 \ALUSHT/ALU/U704  ( .ZN(\ALUSHT/ALU/pkaddinb[6] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[6] ) );
    snl_nor02x1 \ALUSHT/ALU/U846  ( .ZN(\ALUSHT/ALU/n1821 ), .A(
        \ALUSHT/ALU/n1875 ), .B(\ALUSHT/ALU/n1803 ) );
    snl_nor02x1 \ALUSHT/ALU/U498  ( .ZN(\ALUSHT/ALU/pkdecin[16] ), .A(
        \ALUSHT/ALU/n1838 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_and02x1 \ALUSHT/ALU/U508  ( .Z(\ALUSHT/ALU/pkdecin[5] ), .A(
        \pgaluina[5] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_nand02x1 \ALUSHT/ALU/U638  ( .ZN(\ALUSHT/ALU/n2161 ), .A(
        \ALUSHT/ALU/n2162 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nand02x1 \ALUSHT/ALU/U671  ( .ZN(\ALUSHT/ALU/n2211 ), .A(
        \ALUSHT/ALU/n2212 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1041  ( .ZN(\ALUSHT/ALU/n2252 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1906 ) );
    snl_nor02x2 \ALUSHT/ALU/U377  ( .ZN(\ALUSHT/ALU/n2296 ), .A(
        \ALUSHT/ALU/n2093 ), .B(\ALUSHT/ALU/n2082 ) );
    snl_nand04x0 \ALUSHT/ALU/U541  ( .ZN(\ALUSHT/pkaluout[4] ), .A(
        \ALUSHT/ALU/n2018 ), .B(\ALUSHT/ALU/n2019 ), .C(\ALUSHT/ALU/n2020 ), 
        .D(\ALUSHT/ALU/n2021 ) );
    snl_muxi21x1 \ALUSHT/ALU/U933  ( .ZN(\ALUSHT/ALU/n2003 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1891 ) );
    snl_invx05 \ALUSHT/ALU/U566  ( .ZN(\ALUSHT/ALU/n2076 ), .A(\poalufnc[0] )
         );
    snl_nor02x1 \ALUSHT/ALU/U884  ( .ZN(\ALUSHT/ALU/n1865 ), .A(
        \ALUSHT/ALU/n1826 ), .B(\ALUSHT/ALU/inta[25] ) );
    snl_nor02x1 \ALUSHT/ALU/U914  ( .ZN(\ALUSHT/ALU/n1879 ), .A(
        \ALUSHT/ALU/n1878 ), .B(\pgaluina[14] ) );
    snl_nor02x1 \ALUSHT/ALU/U441  ( .ZN(\ALUSHT/ALU/pkaddina[10] ), .A(
        \ALUSHT/ALU/n1843 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U466  ( .ZN(\ALUSHT/ALU/pkincin[17] ), .A(
        \ALUSHT/ALU/n1834 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1837 ), .E(\ALUSHT/ALU/n1873 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai012x1 \ALUSHT/ALU/U656  ( .ZN(\ALUSHT/ALU/n2189 ), .A(
        \ALUSHT/ALU/intb[27] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1008  ( .ZN(\ALUSHT/ALU/n1959 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1871 ) );
    snl_nor04x0 \ALUSHT/ALU/U756  ( .ZN(\ALUSHT/ALU/n2139 ), .A(
        \ALUSHT/ALU/n1847 ), .B(\ALUSHT/ALU/n1848 ), .C(\ALUSHT/ALU/n1849 ), 
        .D(\ALUSHT/ALU/n1850 ) );
    snl_nand02x1 \ALUSHT/ALU/U828  ( .ZN(\ALUSHT/ALU/n2256 ), .A(
        \ALUSHT/ALU/n2060 ), .B(\ALUSHT/ALU/n1854 ) );
    snl_aoi112x0 \ALUSHT/ALU/U814  ( .ZN(\ALUSHT/ALU/n1989 ), .A(
        \ALUSHT/ALU/pkaddsum[12] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2285 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U984  ( .ZN(\ALUSHT/ALU/n2200 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[24] )
         );
    snl_invx05 \ALUSHT/ALU/U833  ( .ZN(\ALUSHT/ALU/n2099 ), .A(
        \ALUSHT/ALU/n2233 ) );
    snl_muxi21x1 \ALUSHT/ALU/U370  ( .ZN(\ALUSHT/ALU/n2022 ), .A(
        \ALUSHT/ALU/n2169 ), .B(\ALUSHT/ALU/n2170 ), .S(\pgaluina[3] ) );
    snl_invx1 \ALUSHT/ALU/U389  ( .ZN(\ALUSHT/ALU/n1803 ), .A(exetype1) );
    snl_aoi012x1 \ALUSHT/ALU/U408  ( .ZN(\ALUSHT/ALU/n1823 ), .A(
        \pgaluinb[28] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_oai222x0 \ALUSHT/ALU/U483  ( .ZN(\ALUSHT/ALU/pkincin[0] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1906 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1853 ), .E(\ALUSHT/ALU/n1907 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nand04x0 \ALUSHT/ALU/U534  ( .ZN(\ALUSHT/pkaluout[11] ), .A(
        \ALUSHT/ALU/n1990 ), .B(\ALUSHT/ALU/n1991 ), .C(\ALUSHT/ALU/n1992 ), 
        .D(\ALUSHT/ALU/n1993 ) );
    snl_aoi112x0 \ALUSHT/ALU/U771  ( .ZN(\ALUSHT/ALU/n2025 ), .A(
        \ALUSHT/ALU/pkaddsum[3] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2264 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U928  ( .ZN(\ALUSHT/ALU/n2150 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1888 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1013  ( .ZN(\ALUSHT/ALU/n1962 ), .A(
        \ALUSHT/ALU/n2219 ), .B(\ALUSHT/ALU/n2220 ), .S(\ALUSHT/ALU/inta[18] )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1034  ( .ZN(\ALUSHT/ALU/n1988 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[12] ) );
    snl_muxi21x1 \ALUSHT/ALU/U946  ( .ZN(\ALUSHT/ALU/n2168 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1898 ) );
    snl_nor02x1 \ALUSHT/ALU/U604  ( .ZN(\ALUSHT/ALU/pkdecin[31] ), .A(
        \ALUSHT/ALU/n1908 ), .B(\ALUSHT/ALU/pkcmpina[31] ) );
    snl_nand12x1 \ALUSHT/ALU/U623  ( .ZN(\ALUSHT/ALU/n2121 ), .A(
        \ALUSHT/ALU/pkaddsum[15] ), .B(\ALUSHT/ALU/pkaddinb[15] ) );
    snl_aoi112x0 \ALUSHT/ALU/U794  ( .ZN(\ALUSHT/ALU/n1953 ), .A(
        \ALUSHT/ALU/pkaddsum[21] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2276 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U961  ( .ZN(\ALUSHT/ALU/n2182 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[2] ) );
    snl_nor02x1 \ALUSHT/ALU/U513  ( .ZN(\ALUSHT/ALU/pkdecin[0] ), .A(
        \ALUSHT/ALU/n1853 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_or04x1 \ALUSHT/ALU/U738  ( .Z(\ALUSHT/ALU/n2131 ), .A(
        \ALUSHT/ALU/inta[22] ), .B(\ALUSHT/ALU/inta[23] ), .C(
        \ALUSHT/ALU/inta[24] ), .D(\ALUSHT/ALU/inta[25] ) );
    snl_nor02x1 \ALUSHT/ALU/U428  ( .ZN(\ALUSHT/ALU/pkaddina[24] ), .A(
        \ALUSHT/ALU/n1810 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U484  ( .ZN(\ALUSHT/ALU/pkdecin[30] ), .A(
        \ALUSHT/ALU/n1802 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand04x0 \ALUSHT/ALU/U514  ( .ZN(\ALUSHT/pkaluout[31] ), .A(
        \ALUSHT/ALU/n1910 ), .B(\ALUSHT/ALU/n1911 ), .C(\ALUSHT/ALU/n1912 ), 
        .D(\ALUSHT/ALU/n1913 ) );
    snl_invx05 \ALUSHT/ALU/U598  ( .ZN(\ALUSHT/ALU/n1906 ), .A(\pgaluinb[0] )
         );
    snl_nand04x0 \ALUSHT/ALU/U533  ( .ZN(\ALUSHT/pkaluout[12] ), .A(
        \ALUSHT/ALU/n1986 ), .B(\ALUSHT/ALU/n1987 ), .C(\ALUSHT/ALU/n1988 ), 
        .D(\ALUSHT/ALU/n1989 ) );
    snl_nand02x1 \ALUSHT/ALU/U603  ( .ZN(\ALUSHT/ALU/n2091 ), .A(
        \pgaluinb[15] ), .B(\pgaluina[15] ) );
    snl_muxi21x1 \ALUSHT/ALU/U624  ( .ZN(\ALUSHT/ALU/n2041 ), .A(
        \ALUSHT/ALU/n2122 ), .B(\ALUSHT/ALU/pkovf32 ), .S(\ALUSHT/ALU/n1803 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U966  ( .ZN(\ALUSHT/ALU/n1918 ), .A(
        \ALUSHT/ALU/n2183 ), .B(\ALUSHT/ALU/n2184 ), .S(\ALUSHT/ALU/inta[29] )
         );
    snl_ao022x1 \ALUSHT/ALU/U793  ( .Z(\ALUSHT/ALU/n2276 ), .A(
        \ALUSHT/ALU/pkdecout[21] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[21] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_nand02x1 \ALUSHT/ALU/U688  ( .ZN(\ALUSHT/ALU/n2236 ), .A(
        \ALUSHT/ALU/n2237 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U718  ( .ZN(\ALUSHT/ALU/pkaddinb[22] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1829 ) );
    snl_muxi21x1 \ALUSHT/ALU/U941  ( .ZN(\ALUSHT/ALU/n2010 ), .A(
        \ALUSHT/ALU/n2160 ), .B(\ALUSHT/ALU/n2161 ), .S(\pgaluina[6] ) );
    snl_nor02x1 \ALUSHT/ALU/U446  ( .ZN(\ALUSHT/ALU/pkaddina[5] ), .A(
        \ALUSHT/ALU/n1848 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_aoi112x0 \ALUSHT/ALU/U776  ( .ZN(\ALUSHT/ALU/n2029 ), .A(
        \ALUSHT/ALU/pkaddsum[2] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2267 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_oai222x0 \ALUSHT/ALU/U461  ( .ZN(\ALUSHT/ALU/pkincin[22] ), .A(
        \ALUSHT/ALU/n1829 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1812 ), .E(\ALUSHT/ALU/n1868 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nor02x1 \ALUSHT/ALU/U834  ( .ZN(\ALUSHT/ALU/n2055 ), .A(
        \ALUSHT/ALU/n2094 ), .B(\ALUSHT/ALU/n2082 ) );
    snl_nand02x1 \ALUSHT/ALU/U651  ( .ZN(\ALUSHT/ALU/n2181 ), .A(
        \ALUSHT/ALU/n2182 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nor04x0 \ALUSHT/ALU/U751  ( .ZN(\ALUSHT/ALU/n2129 ), .A(
        \ALUSHT/ALU/n1802 ), .B(\ALUSHT/ALU/n1805 ), .C(\ALUSHT/ALU/n1806 ), 
        .D(\ALUSHT/ALU/n1807 ) );
    snl_ao022x1 \ALUSHT/ALU/U813  ( .Z(\ALUSHT/ALU/n2285 ), .A(
        \ALUSHT/ALU/pkdecout[12] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[12] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U983  ( .ZN(\ALUSHT/ALU/n1936 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1826 ) );
    snl_invx05 \ALUSHT/ALU/U898  ( .ZN(\ALUSHT/ALU/intb[20] ), .A(
        \ALUSHT/ALU/n1831 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1033  ( .ZN(\ALUSHT/ALU/n1986 ), .A(
        \ALUSHT/ALU/n2241 ), .B(\ALUSHT/ALU/n2242 ), .S(\pgaluina[12] ) );
    snl_invx05 \ALUSHT/ALU/U908  ( .ZN(\ALUSHT/ALU/intb[17] ), .A(
        \ALUSHT/ALU/n1834 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1014  ( .ZN(\ALUSHT/ALU/n1964 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1833 ) );
    snl_oai012x2 \ALUSHT/ALU/U379  ( .ZN(\ALUSHT/ALU/n2145 ), .A(
        \ALUSHT/ALU/n2079 ), .B(\ALUSHT/ALU/n2094 ), .C(\ALUSHT/ALU/n2146 ) );
    snl_invx1 \ALUSHT/ALU/U387  ( .ZN(\ALUSHT/ALU/n1909 ), .A(
        \ALUSHT/ALU/n1908 ) );
    snl_aoi012x1 \ALUSHT/ALU/U395  ( .ZN(\ALUSHT/ALU/n1809 ), .A(
        \pgaluina[25] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nor02x1 \ALUSHT/ALU/U433  ( .ZN(\ALUSHT/ALU/pkaddina[19] ), .A(
        \ALUSHT/ALU/n1815 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai123x0 \ALUSHT/ALU/U546  ( .ZN(\ALUSHT/aluovf ), .A(
        \ALUSHT/ALU/n2038 ), .B(\ALUSHT/ALU/n2039 ), .C(\ALUSHT/ALU/n2040 ), 
        .D(\ALUSHT/ALU/n1836 ), .E(\ALUSHT/ALU/n2041 ), .F(\ALUSHT/ALU/n2042 )
         );
    snl_nand12x1 \ALUSHT/ALU/U561  ( .ZN(\ALUSHT/ALU/n2075 ), .A(
        \ALUSHT/ALU/n1817 ), .B(\ALUSHT/ALU/n2076 ) );
    snl_invx05 \ALUSHT/ALU/U883  ( .ZN(\ALUSHT/ALU/intb[25] ), .A(
        \ALUSHT/ALU/n1826 ) );
    snl_nor02x1 \ALUSHT/ALU/U913  ( .ZN(\ALUSHT/ALU/n1877 ), .A(
        \ALUSHT/ALU/n1875 ), .B(\pgaluina[15] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1028  ( .ZN(\ALUSHT/ALU/n1983 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1881 ) );
    snl_oai012x1 \ALUSHT/ALU/U676  ( .ZN(\ALUSHT/ALU/n2219 ), .A(
        \ALUSHT/ALU/intb[18] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U934  ( .ZN(\ALUSHT/ALU/n2002 ), .A(
        \ALUSHT/ALU/n2154 ), .B(\ALUSHT/ALU/n2155 ), .S(\pgaluina[8] ) );
    snl_nor04x0 \ALUSHT/ALU/U808  ( .ZN(\ALUSHT/ALU/n1977 ), .A(
        \ALUSHT/ALU/n2229 ), .B(\ALUSHT/ALU/n2231 ), .C(\ALUSHT/ALU/n2232 ), 
        .D(\ALUSHT/ALU/n2234 ) );
    snl_muxi21x1 \ALUSHT/ALU/U998  ( .ZN(\ALUSHT/ALU/n1950 ), .A(
        \ALUSHT/ALU/n2207 ), .B(\ALUSHT/ALU/n2208 ), .S(\ALUSHT/ALU/inta[21] )
         );
    snl_invx05 \ALUSHT/ALU/U584  ( .ZN(\ALUSHT/ALU/n1902 ), .A(\pgaluinb[2] )
         );
    snl_oai012x1 \ALUSHT/ALU/U693  ( .ZN(\ALUSHT/ALU/n2244 ), .A(
        \pgaluinb[11] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U703  ( .ZN(\ALUSHT/ALU/pkaddinb[7] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[7] ) );
    snl_nand02x1 \ALUSHT/ALU/U841  ( .ZN(\ALUSHT/ALU/n2119 ), .A(
        \ALUSHT/ALU/n2084 ), .B(\ALUSHT/ALU/n2080 ) );
    snl_muxi21x1 \ALUSHT/ALU/U724  ( .ZN(\ALUSHT/ALU/pkaddinb[17] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\ALUSHT/ALU/intb[17] )
         );
    snl_aoi012x1 \ALUSHT/ALU/U414  ( .ZN(\ALUSHT/ALU/n1829 ), .A(
        \pgaluinb[22] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U421  ( .ZN(\ALUSHT/ALU/pkaddina[31] ), .A(
        \ALUSHT/ALU/pkcmpina[31] ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nand04x0 \ALUSHT/ALU/U528  ( .ZN(\ALUSHT/pkaluout[17] ), .A(
        \ALUSHT/ALU/n1966 ), .B(\ALUSHT/ALU/n1967 ), .C(\ALUSHT/ALU/n1968 ), 
        .D(\ALUSHT/ALU/n1969 ) );
    snl_nor02x1 \ALUSHT/ALU/U866  ( .ZN(\ALUSHT/ALU/n1903 ), .A(
        \ALUSHT/ALU/n1902 ), .B(\pgaluina[2] ) );
    snl_xor2x0 \ALUSHT/ALU/U1046  ( .Z(\ALUSHT/ALU/n2111 ), .A(
        \ALUSHT/ALU/intb[22] ), .B(\ALUSHT/ALU/n1827 ) );
    snl_xor3x1 \ALUSHT/ALU/U618  ( .Z(\ALUSHT/ALU/n2113 ), .A(
        \ALUSHT/ALU/n2114 ), .B(\ALUSHT/ALU/n2115 ), .C(\ALUSHT/ALU/n1900 ) );
    snl_aoi112x0 \ALUSHT/ALU/U788  ( .ZN(\ALUSHT/ALU/n1941 ), .A(
        \ALUSHT/ALU/pkaddsum[24] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2273 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U853  ( .ZN(\ALUSHT/ALU/n1893 ), .A(
        \ALUSHT/ALU/n1892 ), .B(\pgaluina[7] ) );
    snl_muxi21x1 \ALUSHT/ALU/U948  ( .ZN(\ALUSHT/ALU/n2018 ), .A(
        \ALUSHT/ALU/n2166 ), .B(\ALUSHT/ALU/n2167 ), .S(\pgaluina[4] ) );
    snl_xnor2x0 \ALUSHT/ALU/U1054  ( .ZN(\ALUSHT/ALU/n2295 ), .A(
        \ALUSHT/ALU/n1898 ), .B(\ALUSHT/ALU/n1896 ) );
    snl_nand02x1 \ALUSHT/ALU/U681  ( .ZN(\ALUSHT/ALU/n2226 ), .A(
        \ALUSHT/ALU/n2227 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U711  ( .ZN(\ALUSHT/ALU/pkaddinb[29] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1822 ) );
    snl_or04x1 \ALUSHT/ALU/U736  ( .Z(\ALUSHT/ALU/n2040 ), .A(
        \ALUSHT/ALU/n1905 ), .B(\ALUSHT/ALU/n1903 ), .C(\ALUSHT/ALU/n1901 ), 
        .D(\ALUSHT/ALU/n1899 ) );
    snl_invx05 \ALUSHT/ALU/U874  ( .ZN(\ALUSHT/ALU/n2063 ), .A(
        \ALUSHT/ALU/n1862 ) );
    snl_aoi012x1 \ALUSHT/ALU/U406  ( .ZN(\ALUSHT/ALU/n1820 ), .A(
        \pgaluinb[30] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_oai222x0 \ALUSHT/ALU/U468  ( .ZN(\ALUSHT/ALU/pkincin[15] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1875 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1876 ), .E(\ALUSHT/ALU/n1877 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_invx05 \ALUSHT/ALU/U596  ( .ZN(\ALUSHT/ALU/n1886 ), .A(\pgaluinb[10] )
         );
    snl_ao022x1 \ALUSHT/ALU/U758  ( .Z(\ALUSHT/ALU/n2258 ), .A(
        \ALUSHT/ALU/pkdecout[9] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[9] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U554  ( .ZN(\ALUSHT/ALU/pkaddinb[15] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[15] ) );
    snl_invx05 \ALUSHT/ALU/U573  ( .ZN(\ALUSHT/ALU/n1894 ), .A(\pgaluinb[6] )
         );
    snl_oai012x1 \ALUSHT/ALU/U643  ( .ZN(\ALUSHT/ALU/n2169 ), .A(\pgaluinb[3] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_invx05 \ALUSHT/ALU/U891  ( .ZN(\ALUSHT/ALU/inta[22] ), .A(
        \ALUSHT/ALU/n1812 ) );
    snl_invx05 \ALUSHT/ALU/U901  ( .ZN(\ALUSHT/ALU/inta[19] ), .A(
        \ALUSHT/ALU/n1815 ) );
    snl_muxi21x1 \ALUSHT/ALU/U926  ( .ZN(\ALUSHT/ALU/n2137 ), .A(
        \ALUSHT/ALU/n2125 ), .B(\ALUSHT/ALU/n2123 ), .S(exetype1) );
    snl_invx05 \ALUSHT/ALU/U568  ( .ZN(\ALUSHT/ALU/n1845 ), .A(\pgaluina[8] )
         );
    snl_oai012x1 \ALUSHT/ALU/U664  ( .ZN(\ALUSHT/ALU/n2201 ), .A(
        \ALUSHT/ALU/intb[23] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1021  ( .ZN(\ALUSHT/ALU/n1970 ), .A(
        \ALUSHT/ALU/n2225 ), .B(\ALUSHT/ALU/n2226 ), .S(\ALUSHT/ALU/inta[16] )
         );
    snl_oai222x0 \ALUSHT/ALU/U454  ( .ZN(\ALUSHT/ALU/pkincin[29] ), .A(
        \ALUSHT/ALU/n1822 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1805 ), .E(\ALUSHT/ALU/n1861 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai012x1 \ALUSHT/ALU/U658  ( .ZN(\ALUSHT/ALU/n2192 ), .A(
        \ALUSHT/ALU/intb[26] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1006  ( .ZN(\ALUSHT/ALU/n2032 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1904 ) );
    snl_ao022x1 \ALUSHT/ALU/U764  ( .Z(\ALUSHT/ALU/n2261 ), .A(
        \ALUSHT/ALU/pkdecout[6] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[6] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_xor3x1 \ALUSHT/ALU/U826  ( .Z(\ALUSHT/ALU/n2072 ), .A(
        \ALUSHT/ALU/n2113 ), .B(\ALUSHT/ALU/n2293 ), .C(\ALUSHT/ALU/n2295 ) );
    snl_oai222x0 \ALUSHT/ALU/U473  ( .ZN(\ALUSHT/ALU/pkincin[10] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1886 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1843 ), .E(\ALUSHT/ALU/n1887 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_ao022x1 \ALUSHT/ALU/U801  ( .Z(\ALUSHT/ALU/n2280 ), .A(
        \ALUSHT/ALU/pkdecout[18] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[18] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_muxi21x1 \ALUSHT/ALU/U991  ( .ZN(\ALUSHT/ALU/n1944 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1828 ) );
    snl_nor04x0 \ALUSHT/ALU/U743  ( .ZN(\ALUSHT/ALU/n2088 ), .A(
        \ALUSHT/ALU/n1894 ), .B(\ALUSHT/ALU/n1896 ), .C(\ALUSHT/ALU/n1898 ), 
        .D(\ALUSHT/ALU/n1900 ) );
    snl_muxi21x1 \ALUSHT/ALU/U366  ( .ZN(\ALUSHT/ALU/n1990 ), .A(
        \ALUSHT/ALU/n2244 ), .B(\ALUSHT/ALU/n2245 ), .S(\pgaluina[11] ) );
    snl_muxi21x1 \ALUSHT/ALU/U367  ( .ZN(\ALUSHT/ALU/n1994 ), .A(
        \ALUSHT/ALU/n2247 ), .B(\ALUSHT/ALU/n2248 ), .S(\pgaluina[10] ) );
    snl_muxi21x1 \ALUSHT/ALU/U369  ( .ZN(\ALUSHT/ALU/n2014 ), .A(
        \ALUSHT/ALU/n2163 ), .B(\ALUSHT/ALU/n2164 ), .S(\pgaluina[5] ) );
    snl_muxi21x1 \ALUSHT/ALU/U372  ( .ZN(\ALUSHT/ALU/n2030 ), .A(
        \ALUSHT/ALU/n2213 ), .B(\ALUSHT/ALU/n2214 ), .S(\pgaluina[1] ) );
    snl_aoi012x1 \ALUSHT/ALU/U397  ( .ZN(\ALUSHT/ALU/n1811 ), .A(
        \pgaluina[23] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nor02x1 \ALUSHT/ALU/U496  ( .ZN(\ALUSHT/ALU/pkdecin[18] ), .A(
        \ALUSHT/ALU/n1816 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_invx05 \ALUSHT/ALU/U848  ( .ZN(\ALUSHT/ALU/n2080 ), .A(
        \ALUSHT/ALU/n2079 ) );
    snl_muxi21x1 \ALUSHT/ALU/U974  ( .ZN(\ALUSHT/ALU/n1926 ), .A(
        \ALUSHT/ALU/n2189 ), .B(\ALUSHT/ALU/n2190 ), .S(\ALUSHT/ALU/inta[27] )
         );
    snl_and02x1 \ALUSHT/ALU/U506  ( .Z(\ALUSHT/ALU/pkdecin[7] ), .A(
        \pgaluina[7] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_nand04x0 \ALUSHT/ALU/U521  ( .ZN(\ALUSHT/pkaluout[24] ), .A(
        \ALUSHT/ALU/n1938 ), .B(\ALUSHT/ALU/n1939 ), .C(\ALUSHT/ALU/n1940 ), 
        .D(\ALUSHT/ALU/n1941 ) );
    snl_and02x1 \ALUSHT/ALU/U611  ( .Z(\ALUSHT/ALU/n2097 ), .A(
        \ALUSHT/ALU/n2098 ), .B(\ALUSHT/ALU/n2099 ) );
    snl_nand02x1 \ALUSHT/ALU/U636  ( .ZN(\ALUSHT/ALU/n2158 ), .A(
        \ALUSHT/ALU/n2159 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_ao022x1 \ALUSHT/ALU/U781  ( .Z(\ALUSHT/ALU/n2270 ), .A(
        \ALUSHT/ALU/pkdecout[27] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[27] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_mux21x1 \ALUSHT/ALU/U953  ( .Z(\ALUSHT/ALU/n2176 ), .A(
        \ALUSHT/ALU/n2148 ), .B(\ALUSHT/ALU/n2228 ), .S(\ALUSHT/ALU/n1854 ) );
    snl_invx05 \ALUSHT/ALU/U586  ( .ZN(\ALUSHT/ALU/n1904 ), .A(\pgaluinb[1] )
         );
    snl_muxi21x1 \ALUSHT/ALU/U726  ( .ZN(\ALUSHT/ALU/pkaddinb[14] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1878 ) );
    snl_muxi21x1 \ALUSHT/ALU/U958  ( .ZN(\ALUSHT/ALU/n1915 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1859 ) );
    snl_xor2x0 \ALUSHT/ALU/U1044  ( .Z(\ALUSHT/ALU/n2107 ), .A(
        \ALUSHT/ALU/intb[30] ), .B(\ALUSHT/ALU/pkcmpinb[31] ) );
    snl_nor02x1 \ALUSHT/ALU/U864  ( .ZN(\ALUSHT/ALU/n1859 ), .A(
        \ALUSHT/ALU/n1820 ), .B(\ALUSHT/ALU/inta[30] ) );
    snl_aoi012x1 \ALUSHT/ALU/U416  ( .ZN(\ALUSHT/ALU/n1831 ), .A(
        \pgaluinb[20] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U431  ( .ZN(\ALUSHT/ALU/pkaddina[21] ), .A(
        \ALUSHT/ALU/n1813 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U843  ( .ZN(\ALUSHT/ALU/pkaddina[15] ), .A(
        \ALUSHT/ALU/n1836 ), .B(\ALUSHT/ALU/n1876 ) );
    snl_oai222x0 \ALUSHT/ALU/U478  ( .ZN(\ALUSHT/ALU/pkincin[5] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1896 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1848 ), .E(\ALUSHT/ALU/n1897 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai012x1 \ALUSHT/ALU/U691  ( .ZN(\ALUSHT/ALU/n2241 ), .A(
        \pgaluinb[12] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U701  ( .ZN(\ALUSHT/ALU/pkaddinb[9] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[9] ) );
    snl_nor04x0 \ALUSHT/ALU/U748  ( .ZN(\ALUSHT/ALU/n2052 ), .A(
        \ALUSHT/ALU/n2257 ), .B(\ALUSHT/ALU/n2255 ), .C(\ALUSHT/ALU/n1823 ), 
        .D(\ALUSHT/ALU/n1824 ) );
    snl_nand04x0 \ALUSHT/ALU/U544  ( .ZN(\ALUSHT/pkaluout[1] ), .A(
        \ALUSHT/ALU/n2030 ), .B(\ALUSHT/ALU/n2031 ), .C(\ALUSHT/ALU/n2032 ), 
        .D(\ALUSHT/ALU/n2033 ) );
    snl_muxi21x1 \ALUSHT/ALU/U936  ( .ZN(\ALUSHT/ALU/n2159 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[7] ) );
    snl_nand02x1 \ALUSHT/ALU/U653  ( .ZN(\ALUSHT/ALU/n2184 ), .A(
        \ALUSHT/ALU/n2185 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_oai012x1 \ALUSHT/ALU/U674  ( .ZN(\ALUSHT/ALU/n2216 ), .A(
        \ALUSHT/ALU/intb[19] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_nor02x1 \ALUSHT/ALU/U881  ( .ZN(\ALUSHT/ALU/n1864 ), .A(
        \ALUSHT/ALU/n1825 ), .B(\ALUSHT/ALU/inta[26] ) );
    snl_invx05 \ALUSHT/ALU/U911  ( .ZN(\ALUSHT/ALU/intb[16] ), .A(
        \ALUSHT/ALU/n1835 ) );
    snl_nand02x1 \ALUSHT/ALU/U563  ( .ZN(\ALUSHT/ALU/n2048 ), .A(
        \ALUSHT/ALU/n1817 ), .B(\ALUSHT/ALU/n2076 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1016  ( .ZN(\ALUSHT/ALU/n1967 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1873 ) );
    snl_nand02x2 \ALUSHT/ALU/U382  ( .ZN(\ALUSHT/ALU/n1818 ), .A(
        \ALUSHT/ALU/n2084 ), .B(\ALUSHT/ALU/n2076 ) );
    snl_nor02x2 \ALUSHT/ALU/U385  ( .ZN(\ALUSHT/ALU/n1974 ), .A(
        \ALUSHT/ALU/n2093 ), .B(\ALUSHT/ALU/n2048 ) );
    snl_nor02x1 \ALUSHT/ALU/U438  ( .ZN(\ALUSHT/ALU/pkaddina[13] ), .A(
        \ALUSHT/ALU/n1840 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U444  ( .ZN(\ALUSHT/ALU/pkaddina[7] ), .A(
        \ALUSHT/ALU/n1846 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U463  ( .ZN(\ALUSHT/ALU/pkincin[20] ), .A(
        \ALUSHT/ALU/n1831 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1814 ), .E(\ALUSHT/ALU/n1870 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_invx05 \ALUSHT/ALU/U578  ( .ZN(\ALUSHT/ALU/n1850 ), .A(\pgaluina[3] )
         );
    snl_oai012x1 \ALUSHT/ALU/U648  ( .ZN(\ALUSHT/ALU/n2177 ), .A(
        \ALUSHT/ALU/intb[30] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_ao022x1 \ALUSHT/ALU/U811  ( .Z(\ALUSHT/ALU/n2284 ), .A(
        \ALUSHT/ALU/pkdecout[13] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[13] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1031  ( .ZN(\ALUSHT/ALU/n2243 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1882 ) );
    snl_muxi21x1 \ALUSHT/ALU/U981  ( .ZN(\ALUSHT/ALU/n1935 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1865 ) );
    snl_nor04x0 \ALUSHT/ALU/U753  ( .ZN(\ALUSHT/ALU/n2127 ), .A(
        \ALUSHT/ALU/n1814 ), .B(\ALUSHT/ALU/n1812 ), .C(\ALUSHT/ALU/n1813 ), 
        .D(\ALUSHT/ALU/n1815 ) );
    snl_ao022x1 \ALUSHT/ALU/U774  ( .Z(\ALUSHT/ALU/n2266 ), .A(
        \ALUSHT/ALU/pkdecout[30] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[30] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_invx05 \ALUSHT/ALU/U836  ( .ZN(\ALUSHT/ALU/n2146 ), .A(
        \ALUSHT/ALU/n2095 ) );
    snl_nor02x1 \ALUSHT/ALU/U486  ( .ZN(\ALUSHT/ALU/pkdecin[28] ), .A(
        \ALUSHT/ALU/n1806 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand04x0 \ALUSHT/ALU/U516  ( .ZN(\ALUSHT/pkaluout[29] ), .A(
        \ALUSHT/ALU/n1918 ), .B(\ALUSHT/ALU/n1919 ), .C(\ALUSHT/ALU/n1920 ), 
        .D(\ALUSHT/ALU/n1921 ) );
    snl_nand04x0 \ALUSHT/ALU/U531  ( .ZN(\ALUSHT/pkaluout[14] ), .A(
        \ALUSHT/ALU/n1978 ), .B(\ALUSHT/ALU/n1979 ), .C(\ALUSHT/ALU/n1980 ), 
        .D(\ALUSHT/ALU/n1981 ) );
    snl_nand04x0 \ALUSHT/ALU/U601  ( .ZN(\ALUSHT/ALU/n2085 ), .A(
        \ALUSHT/ALU/n2086 ), .B(\ALUSHT/ALU/n2087 ), .C(\ALUSHT/ALU/n2088 ), 
        .D(\ALUSHT/ALU/n2089 ) );
    snl_ao022x1 \ALUSHT/ALU/U791  ( .Z(\ALUSHT/ALU/n2275 ), .A(
        \ALUSHT/ALU/pkdecout[22] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[22] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_invx05 \ALUSHT/ALU/U858  ( .ZN(\ALUSHT/ALU/n1854 ), .A(
        \ALUSHT/ALU/pkcmpina[31] ) );
    snl_muxi21x1 \ALUSHT/ALU/U943  ( .ZN(\ALUSHT/ALU/n2165 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[5] ) );
    snl_muxi21x1 \ALUSHT/ALU/U964  ( .ZN(\ALUSHT/ALU/n2185 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1822 ) );
    snl_nor02x1 \ALUSHT/ALU/U494  ( .ZN(\ALUSHT/ALU/pkdecin[20] ), .A(
        \ALUSHT/ALU/n1814 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand04x0 \ALUSHT/ALU/U523  ( .ZN(\ALUSHT/pkaluout[22] ), .A(
        \ALUSHT/ALU/n1946 ), .B(\ALUSHT/ALU/n1947 ), .C(\ALUSHT/ALU/n1948 ), 
        .D(\ALUSHT/ALU/n1949 ) );
    snl_and02x1 \ALUSHT/ALU/U613  ( .Z(\ALUSHT/ALU/n2102 ), .A(
        \ALUSHT/ALU/n2103 ), .B(\ALUSHT/ALU/n1803 ) );
    snl_nand04x0 \ALUSHT/ALU/U626  ( .ZN(\ALUSHT/ALU/n2125 ), .A(
        \ALUSHT/ALU/n2126 ), .B(\ALUSHT/ALU/n2127 ), .C(\ALUSHT/ALU/n2128 ), 
        .D(\ALUSHT/ALU/n2129 ) );
    snl_ao022x1 \ALUSHT/ALU/U783  ( .Z(\ALUSHT/ALU/n2271 ), .A(
        \ALUSHT/ALU/pkdecout[26] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[26] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_muxi21x1 \ALUSHT/ALU/U951  ( .ZN(\ALUSHT/ALU/n2023 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1901 ) );
    snl_nor02x1 \ALUSHT/ALU/U504  ( .ZN(\ALUSHT/ALU/pkdecin[9] ), .A(
        \ALUSHT/ALU/n1844 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand02x1 \ALUSHT/ALU/U634  ( .ZN(\ALUSHT/ALU/n2155 ), .A(
        \ALUSHT/ALU/n2156 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U976  ( .ZN(\ALUSHT/ALU/n2194 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[26] )
         );
    snl_nand02x1 \ALUSHT/ALU/U698  ( .ZN(\ALUSHT/ALU/n2251 ), .A(
        \ALUSHT/ALU/n2252 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U708  ( .ZN(\ALUSHT/ALU/pkaddinb[31] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\ALUSHT/ALU/n2060 ) );
    snl_oai222x0 \ALUSHT/ALU/U456  ( .ZN(\ALUSHT/ALU/pkincin[27] ), .A(
        \ALUSHT/ALU/n1824 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1807 ), .E(\ALUSHT/ALU/n1863 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai222x0 \ALUSHT/ALU/U471  ( .ZN(\ALUSHT/ALU/pkincin[12] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1882 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1841 ), .E(\ALUSHT/ALU/n1883 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_and08x1 \ALUSHT/ALU/U741  ( .Z(\ALUSHT/ALU/n2142 ), .A(
        \ALUSHT/ALU/n1847 ), .B(\ALUSHT/ALU/n1846 ), .C(\ALUSHT/ALU/n1845 ), 
        .D(\ALUSHT/ALU/n1844 ), .E(\ALUSHT/ALU/n1843 ), .F(\ALUSHT/ALU/n1842 ), 
        .G(\ALUSHT/ALU/n1841 ), .H(\ALUSHT/ALU/n1840 ) );
    snl_ao022x1 \ALUSHT/ALU/U803  ( .Z(\ALUSHT/ALU/n2281 ), .A(
        \ALUSHT/ALU/pkdecout[17] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[17] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_muxi21x1 \ALUSHT/ALU/U993  ( .ZN(\ALUSHT/ALU/n1947 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1868 ) );
    snl_ao022x1 \ALUSHT/ALU/U766  ( .Z(\ALUSHT/ALU/n2262 ), .A(
        \ALUSHT/ALU/pkdecout[5] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[5] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_xnor2x0 \ALUSHT/ALU/U556  ( .ZN(\ALUSHT/ALU/n2068 ), .A(
        \ALUSHT/ALU/pkeqflg ), .B(\poalufnc[0] ) );
    snl_xor3x1 \ALUSHT/ALU/U824  ( .Z(\ALUSHT/ALU/n2293 ), .A(
        \ALUSHT/ALU/n2106 ), .B(\ALUSHT/ALU/n2291 ), .C(\ALUSHT/ALU/n2290 ) );
    snl_invx05 \ALUSHT/ALU/U888  ( .ZN(\ALUSHT/ALU/inta[23] ), .A(
        \ALUSHT/ALU/n1811 ) );
    snl_nor02x1 \ALUSHT/ALU/U918  ( .ZN(\ALUSHT/ALU/n1887 ), .A(
        \ALUSHT/ALU/n1886 ), .B(\pgaluina[10] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1004  ( .ZN(\ALUSHT/ALU/n2215 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[1] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1023  ( .ZN(\ALUSHT/ALU/n2237 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[14] ) );
    snl_invx05 \ALUSHT/ALU/U571  ( .ZN(\ALUSHT/ALU/n1892 ), .A(\pgaluinb[7] )
         );
    snl_oai012x1 \ALUSHT/ALU/U641  ( .ZN(\ALUSHT/ALU/n2166 ), .A(\pgaluinb[4] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_oai012x1 \ALUSHT/ALU/U666  ( .ZN(\ALUSHT/ALU/n2204 ), .A(
        \ALUSHT/ALU/intb[22] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_mux21x1 \ALUSHT/ALU/U924  ( .Z(\ALUSHT/ALU/n1856 ), .A(
        \ALUSHT/ALU/n1860 ), .B(\ALUSHT/ALU/n1857 ), .S(\ALUSHT/ALU/n2060 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1038  ( .ZN(\ALUSHT/ALU/n2249 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\pgaluinb[10] ) );
    snl_nor04x0 \ALUSHT/ALU/U734  ( .ZN(\ALUSHT/ALU/n2065 ), .A(
        \ALUSHT/ALU/n1872 ), .B(\ALUSHT/ALU/n1873 ), .C(\ALUSHT/ALU/n1874 ), 
        .D(\ALUSHT/ALU/n1854 ) );
    snl_aoi112x0 \ALUSHT/ALU/U818  ( .ZN(\ALUSHT/ALU/n1997 ), .A(
        \ALUSHT/ALU/pkaddsum[10] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2287 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U893  ( .ZN(\ALUSHT/ALU/n1868 ), .A(
        \ALUSHT/ALU/n1829 ), .B(\ALUSHT/ALU/inta[22] ) );
    snl_nor02x1 \ALUSHT/ALU/U903  ( .ZN(\ALUSHT/ALU/n1871 ), .A(
        \ALUSHT/ALU/n1832 ), .B(\ALUSHT/ALU/inta[19] ) );
    snl_muxi21x1 \ALUSHT/ALU/U988  ( .ZN(\ALUSHT/ALU/n2203 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[23] )
         );
    snl_ao012x1 \ALUSHT/ALU/U403  ( .Z(\ALUSHT/ALU/inta[17] ), .A(
        \pgaluina[17] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_ao012x1 \ALUSHT/ALU/U404  ( .Z(\ALUSHT/ALU/inta[16] ), .A(
        \pgaluina[16] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nor02x1 \ALUSHT/ALU/U423  ( .ZN(\ALUSHT/ALU/pkaddina[29] ), .A(
        \ALUSHT/ALU/n1805 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_invx05 \ALUSHT/ALU/U594  ( .ZN(\ALUSHT/ALU/n1884 ), .A(\pgaluinb[11] )
         );
    snl_invx05 \ALUSHT/ALU/U876  ( .ZN(\ALUSHT/ALU/intb[27] ), .A(
        \ALUSHT/ALU/n1824 ) );
    snl_nor02x1 \ALUSHT/ALU/U424  ( .ZN(\ALUSHT/ALU/pkaddina[28] ), .A(
        \ALUSHT/ALU/n1806 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nand04x0 \ALUSHT/ALU/U538  ( .ZN(\ALUSHT/pkaluout[7] ), .A(
        \ALUSHT/ALU/n2006 ), .B(\ALUSHT/ALU/n2007 ), .C(\ALUSHT/ALU/n2008 ), 
        .D(\ALUSHT/ALU/n2009 ) );
    snl_muxi21x1 \ALUSHT/ALU/U683  ( .ZN(\ALUSHT/ALU/n2229 ), .A(
        \ALUSHT/ALU/n2054 ), .B(\ALUSHT/ALU/n2230 ), .S(\pgaluinb[15] ) );
    snl_nor02x1 \ALUSHT/ALU/U851  ( .ZN(\ALUSHT/ALU/n1889 ), .A(
        \ALUSHT/ALU/n1888 ), .B(\pgaluina[9] ) );
    snl_muxi21x1 \ALUSHT/ALU/U713  ( .ZN(\ALUSHT/ALU/pkaddinb[27] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\ALUSHT/ALU/intb[27] )
         );
    snl_nand02x1 \ALUSHT/ALU/U608  ( .ZN(\ALUSHT/ALU/n2094 ), .A(
        \ALUSHT/ALU/n2074 ), .B(\ALUSHT/ALU/n2044 ) );
    snl_muxi21x1 \ALUSHT/ALU/U684  ( .ZN(\ALUSHT/ALU/n2231 ), .A(
        \ALUSHT/ALU/n2098 ), .B(\ALUSHT/ALU/n2100 ), .S(\pgaluina[15] ) );
    snl_muxi21x1 \ALUSHT/ALU/U714  ( .ZN(\ALUSHT/ALU/pkaddinb[26] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1825 ) );
    snl_aoi112x0 \ALUSHT/ALU/U798  ( .ZN(\ALUSHT/ALU/n2033 ), .A(
        \ALUSHT/ALU/pkaddsum[1] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2278 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U856  ( .ZN(\ALUSHT/ALU/n1899 ), .A(
        \ALUSHT/ALU/n1898 ), .B(\pgaluina[4] ) );
    snl_invx05 \ALUSHT/ALU/U593  ( .ZN(\ALUSHT/ALU/n1842 ), .A(\pgaluina[11] )
         );
    snl_invx05 \ALUSHT/ALU/U871  ( .ZN(\ALUSHT/ALU/inta[28] ), .A(
        \ALUSHT/ALU/n1806 ) );
    snl_nor02x1 \ALUSHT/ALU/U488  ( .ZN(\ALUSHT/ALU/pkdecin[26] ), .A(
        \ALUSHT/ALU/n1808 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand04x0 \ALUSHT/ALU/U518  ( .ZN(\ALUSHT/pkaluout[27] ), .A(
        \ALUSHT/ALU/n1926 ), .B(\ALUSHT/ALU/n1927 ), .C(\ALUSHT/ALU/n1928 ), 
        .D(\ALUSHT/ALU/n1929 ) );
    snl_nor04x0 \ALUSHT/ALU/U733  ( .ZN(\ALUSHT/ALU/n2066 ), .A(
        \ALUSHT/ALU/n1868 ), .B(\ALUSHT/ALU/n1869 ), .C(\ALUSHT/ALU/n1870 ), 
        .D(\ALUSHT/ALU/n1871 ) );
    snl_xnor2x0 \ALUSHT/ALU/U1051  ( .ZN(\ALUSHT/ALU/n2110 ), .A(
        \ALUSHT/ALU/n1888 ), .B(\ALUSHT/ALU/n1884 ) );
    snl_nand02x1 \ALUSHT/ALU/U628  ( .ZN(\ALUSHT/ALU/n2134 ), .A(
        \ALUSHT/ALU/n1909 ), .B(\pgaluina[15] ) );
    snl_invx05 \ALUSHT/ALU/U894  ( .ZN(\ALUSHT/ALU/inta[21] ), .A(
        \ALUSHT/ALU/n1813 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1018  ( .ZN(\ALUSHT/ALU/n1968 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1834 ) );
    snl_invx05 \ALUSHT/ALU/U904  ( .ZN(\ALUSHT/ALU/inta[18] ), .A(
        \ALUSHT/ALU/n1816 ) );
    snl_nand02x2 \ALUSHT/ALU/U375  ( .ZN(\ALUSHT/ALU/n1908 ), .A(
        \ALUSHT/ALU/n2083 ), .B(\ALUSHT/ALU/n2077 ) );
    snl_aoi012x1 \ALUSHT/ALU/U399  ( .ZN(\ALUSHT/ALU/n1813 ), .A(
        \pgaluina[21] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U418  ( .ZN(\ALUSHT/ALU/n1833 ), .A(
        \pgaluinb[18] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U451  ( .ZN(\ALUSHT/ALU/pkaddina[0] ), .A(
        \ALUSHT/ALU/n1853 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U551  ( .ZN(\ALUSHT/ALU/n2057 ), .A(
        \ALUSHT/ALU/pkeqflg ), .B(\ALUSHT/ALU/pkgtflg ) );
    snl_invx05 \ALUSHT/ALU/U576  ( .ZN(\ALUSHT/ALU/n1849 ), .A(\pgaluina[4] )
         );
    snl_nand02x1 \ALUSHT/ALU/U646  ( .ZN(\ALUSHT/ALU/n2173 ), .A(
        \ALUSHT/ALU/n2100 ), .B(\ALUSHT/ALU/n2174 ) );
    snl_nand02x1 \ALUSHT/ALU/U661  ( .ZN(\ALUSHT/ALU/n2196 ), .A(
        \ALUSHT/ALU/n2197 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_xor2x0 \ALUSHT/ALU/U923  ( .Z(\ALUSHT/ALU/n2254 ), .A(
        \ALUSHT/ALU/n2076 ), .B(\ALUSHT/ALU/n2253 ) );
    snl_xor2x0 \ALUSHT/ALU/U823  ( .Z(\ALUSHT/ALU/n2291 ), .A(
        \ALUSHT/ALU/n2289 ), .B(\ALUSHT/ALU/n2292 ) );
    snl_invx05 \ALUSHT/ALU/U838  ( .ZN(\ALUSHT/ALU/n2174 ), .A(
        \ALUSHT/ALU/n2296 ) );
    snl_oai222x0 \ALUSHT/ALU/U476  ( .ZN(\ALUSHT/ALU/pkincin[7] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1892 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1846 ), .E(\ALUSHT/ALU/n1893 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nand03x0 \ALUSHT/ALU/U746  ( .ZN(\ALUSHT/ALU/n2255 ), .A(
        \ALUSHT/ALU/intb[30] ), .B(\ALUSHT/ALU/n2256 ), .C(
        \ALUSHT/ALU/intb[29] ) );
    snl_aoi112x0 \ALUSHT/ALU/U761  ( .ZN(\ALUSHT/ALU/n2005 ), .A(
        \ALUSHT/ALU/pkaddsum[8] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2259 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_aoi112x0 \ALUSHT/ALU/U804  ( .ZN(\ALUSHT/ALU/n1969 ), .A(
        \ALUSHT/ALU/pkaddsum[17] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2281 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U994  ( .ZN(\ALUSHT/ALU/n1946 ), .A(
        \ALUSHT/ALU/n2204 ), .B(\ALUSHT/ALU/n2205 ), .S(\ALUSHT/ALU/inta[22] )
         );
    snl_nor02x1 \ALUSHT/ALU/U493  ( .ZN(\ALUSHT/ALU/pkdecin[21] ), .A(
        \ALUSHT/ALU/n1813 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nor02x1 \ALUSHT/ALU/U503  ( .ZN(\ALUSHT/ALU/pkdecin[10] ), .A(
        \ALUSHT/ALU/n1843 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_oai012x1 \ALUSHT/ALU/U633  ( .ZN(\ALUSHT/ALU/n2154 ), .A(\pgaluinb[8] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U938  ( .ZN(\ALUSHT/ALU/n2008 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[7] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1003  ( .ZN(\ALUSHT/ALU/n1956 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1831 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1024  ( .ZN(\ALUSHT/ALU/n1979 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1879 ) );
    snl_muxi21x1 \ALUSHT/ALU/U971  ( .ZN(\ALUSHT/ALU/n1924 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1823 ) );
    snl_nand04x0 \ALUSHT/ALU/U524  ( .ZN(\ALUSHT/pkaluout[21] ), .A(
        \ALUSHT/ALU/n1950 ), .B(\ALUSHT/ALU/n1951 ), .C(\ALUSHT/ALU/n1952 ), 
        .D(\ALUSHT/ALU/n1953 ) );
    snl_muxi21x1 \ALUSHT/ALU/U956  ( .ZN(\ALUSHT/ALU/n1912 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2175 ), .S(
        \ALUSHT/ALU/pkcmpinb[31] ) );
    snl_invx05 \ALUSHT/ALU/U588  ( .ZN(\ALUSHT/ALU/n1878 ), .A(\pgaluinb[14] )
         );
    snl_and02x1 \ALUSHT/ALU/U614  ( .Z(\ALUSHT/ALU/n2104 ), .A(
        \ALUSHT/ALU/n1855 ), .B(\ALUSHT/ALU/n1803 ) );
    snl_aoi112x0 \ALUSHT/ALU/U784  ( .ZN(\ALUSHT/ALU/n1933 ), .A(
        \ALUSHT/ALU/pkaddsum[26] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2271 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U728  ( .ZN(\ALUSHT/ALU/pkaddinb[12] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[12] ) );
    snl_nor02x1 \ALUSHT/ALU/U443  ( .ZN(\ALUSHT/ALU/pkaddina[8] ), .A(
        \ALUSHT/ALU/n1845 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U481  ( .ZN(\ALUSHT/ALU/pkincin[2] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1902 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1851 ), .E(\ALUSHT/ALU/n1903 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_and02x1 \ALUSHT/ALU/U621  ( .Z(\ALUSHT/ALU/n2069 ), .A(
        \ALUSHT/ALU/n1819 ), .B(\ALUSHT/ALU/n2119 ) );
    snl_invx05 \ALUSHT/ALU/U878  ( .ZN(\ALUSHT/ALU/n2062 ), .A(
        \ALUSHT/ALU/n1863 ) );
    snl_and02x1 \ALUSHT/ALU/U511  ( .Z(\ALUSHT/ALU/pkdecin[2] ), .A(
        \pgaluina[2] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_nand04x0 \ALUSHT/ALU/U536  ( .ZN(\ALUSHT/pkaluout[9] ), .A(
        \ALUSHT/ALU/n1998 ), .B(\ALUSHT/ALU/n1999 ), .C(\ALUSHT/ALU/n2000 ), 
        .D(\ALUSHT/ALU/n2001 ) );
    snl_muxi21x1 \ALUSHT/ALU/U963  ( .ZN(\ALUSHT/ALU/n2028 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[2] ) );
    snl_nor02x1 \ALUSHT/ALU/U558  ( .ZN(\ALUSHT/ALU/n2074 ), .A(
        \ALUSHT/ALU/n2073 ), .B(\poalufnc[3] ) );
    snl_and02x1 \ALUSHT/ALU/U606  ( .Z(\ALUSHT/ALU/n2092 ), .A(\poalufnc[3] ), 
        .B(\ALUSHT/ALU/n2044 ) );
    snl_muxi21x1 \ALUSHT/ALU/U944  ( .ZN(\ALUSHT/ALU/n2015 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1897 ) );
    snl_aoi112x0 \ALUSHT/ALU/U796  ( .ZN(\ALUSHT/ALU/n1957 ), .A(
        \ALUSHT/ALU/pkaddsum[20] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2277 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_oai012x1 \ALUSHT/ALU/U668  ( .ZN(\ALUSHT/ALU/n2207 ), .A(
        \ALUSHT/ALU/intb[21] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1036  ( .ZN(\ALUSHT/ALU/n1991 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1885 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1011  ( .ZN(\ALUSHT/ALU/n2221 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[18] )
         );
    snl_oai222x0 \ALUSHT/ALU/U458  ( .ZN(\ALUSHT/ALU/pkincin[25] ), .A(
        \ALUSHT/ALU/n1826 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1809 ), .E(\ALUSHT/ALU/n1865 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai222x0 \ALUSHT/ALU/U464  ( .ZN(\ALUSHT/ALU/pkincin[19] ), .A(
        \ALUSHT/ALU/n1832 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1815 ), .E(\ALUSHT/ALU/n1871 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nor04x0 \ALUSHT/ALU/U754  ( .ZN(\ALUSHT/ALU/n2126 ), .A(
        \ALUSHT/ALU/n1816 ), .B(\ALUSHT/ALU/n1837 ), .C(\ALUSHT/ALU/n1838 ), 
        .D(\ALUSHT/ALU/n2049 ) );
    snl_aoi112x0 \ALUSHT/ALU/U773  ( .ZN(\ALUSHT/ALU/n1913 ), .A(
        \ALUSHT/ALU/pkaddsum[31] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2265 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nand02x1 \ALUSHT/ALU/U831  ( .ZN(\ALUSHT/ALU/n2098 ), .A(
        \ALUSHT/ALU/n2096 ), .B(\ALUSHT/ALU/n2090 ) );
    snl_ao022x1 \ALUSHT/ALU/U768  ( .Z(\ALUSHT/ALU/n2263 ), .A(
        \ALUSHT/ALU/pkdecout[4] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[4] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_aoi112x0 \ALUSHT/ALU/U816  ( .ZN(\ALUSHT/ALU/n1993 ), .A(
        \ALUSHT/ALU/pkaddsum[11] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2286 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U986  ( .ZN(\ALUSHT/ALU/n1938 ), .A(
        \ALUSHT/ALU/n2198 ), .B(\ALUSHT/ALU/n2199 ), .S(\ALUSHT/ALU/inta[24] )
         );
    snl_invx05 \ALUSHT/ALU/U564  ( .ZN(\ALUSHT/ALU/n1844 ), .A(\pgaluina[9] )
         );
    snl_aoi012x1 \ALUSHT/ALU/U390  ( .ZN(\ALUSHT/ALU/n1802 ), .A(
        \pgaluina[30] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U411  ( .ZN(\ALUSHT/ALU/n1826 ), .A(
        \pgaluinb[25] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U436  ( .ZN(\ALUSHT/ALU/pkaddina[16] ), .A(
        \ALUSHT/ALU/n1838 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nand04x0 \ALUSHT/ALU/U543  ( .ZN(\ALUSHT/pkaluout[2] ), .A(
        \ALUSHT/ALU/n2026 ), .B(\ALUSHT/ALU/n2027 ), .C(\ALUSHT/ALU/n2028 ), 
        .D(\ALUSHT/ALU/n2029 ) );
    snl_oai012x1 \ALUSHT/ALU/U654  ( .ZN(\ALUSHT/ALU/n2186 ), .A(
        \ALUSHT/ALU/intb[28] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_invx05 \ALUSHT/ALU/U886  ( .ZN(\ALUSHT/ALU/intb[24] ), .A(
        \ALUSHT/ALU/n1827 ) );
    snl_nor02x1 \ALUSHT/ALU/U916  ( .ZN(\ALUSHT/ALU/n1883 ), .A(
        \ALUSHT/ALU/n1882 ), .B(\pgaluina[12] ) );
    snl_nand02x1 \ALUSHT/ALU/U673  ( .ZN(\ALUSHT/ALU/n2214 ), .A(
        \ALUSHT/ALU/n2215 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nand02x1 \ALUSHT/ALU/U696  ( .ZN(\ALUSHT/ALU/n2248 ), .A(
        \ALUSHT/ALU/n2249 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U931  ( .ZN(\ALUSHT/ALU/n2000 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[9] ) );
    snl_muxi21x1 \ALUSHT/ALU/U978  ( .ZN(\ALUSHT/ALU/n1930 ), .A(
        \ALUSHT/ALU/n2192 ), .B(\ALUSHT/ALU/n2193 ), .S(\ALUSHT/ALU/inta[26] )
         );
    snl_muxi21x1 \ALUSHT/ALU/U1043  ( .ZN(\ALUSHT/ALU/n2036 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[0] ) );
    snl_muxi21x1 \ALUSHT/ALU/U706  ( .ZN(\ALUSHT/ALU/pkaddinb[4] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[4] ) );
    snl_invx05 \ALUSHT/ALU/U844  ( .ZN(\ALUSHT/ALU/pkdecin[15] ), .A(
        \ALUSHT/ALU/n2134 ) );
    snl_aoi012x1 \ALUSHT/ALU/U398  ( .ZN(\ALUSHT/ALU/n1812 ), .A(
        \pgaluina[22] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nor02x1 \ALUSHT/ALU/U492  ( .ZN(\ALUSHT/ALU/pkdecin[22] ), .A(
        \ALUSHT/ALU/n1812 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_and02x1 \ALUSHT/ALU/U581  ( .Z(\ALUSHT/ALU/n1858 ), .A(
        \ALUSHT/ALU/n2081 ), .B(\ALUSHT/ALU/n1857 ) );
    snl_nand02x1 \ALUSHT/ALU/U632  ( .ZN(\ALUSHT/ALU/n2149 ), .A(
        \ALUSHT/ALU/n2150 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U721  ( .ZN(\ALUSHT/ALU/pkaddinb[1] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1904 ) );
    snl_invx05 \ALUSHT/ALU/U863  ( .ZN(\ALUSHT/ALU/intb[30] ), .A(
        \ALUSHT/ALU/n1820 ) );
    snl_muxi21x1 \ALUSHT/ALU/U970  ( .ZN(\ALUSHT/ALU/n1922 ), .A(
        \ALUSHT/ALU/n2186 ), .B(\ALUSHT/ALU/n2187 ), .S(\ALUSHT/ALU/inta[28] )
         );
    snl_nor02x1 \ALUSHT/ALU/U502  ( .ZN(\ALUSHT/ALU/pkdecin[11] ), .A(
        \ALUSHT/ALU/n1842 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand04x0 \ALUSHT/ALU/U525  ( .ZN(\ALUSHT/pkaluout[20] ), .A(
        \ALUSHT/ALU/n1954 ), .B(\ALUSHT/ALU/n1955 ), .C(\ALUSHT/ALU/n1956 ), 
        .D(\ALUSHT/ALU/n1957 ) );
    snl_muxi21x1 \ALUSHT/ALU/U957  ( .ZN(\ALUSHT/ALU/n2179 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1820 ) );
    snl_nor02x1 \ALUSHT/ALU/U615  ( .ZN(\ALUSHT/ALU/n2105 ), .A(
        \ALUSHT/ALU/n1908 ), .B(exetype1) );
    snl_muxi21x1 \ALUSHT/ALU/U729  ( .ZN(\ALUSHT/ALU/pkaddinb[11] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[11] ) );
    snl_ao022x1 \ALUSHT/ALU/U785  ( .Z(\ALUSHT/ALU/n2272 ), .A(
        \ALUSHT/ALU/pkdecout[25] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[25] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_aoi012x1 \ALUSHT/ALU/U419  ( .ZN(\ALUSHT/ALU/n1834 ), .A(
        \pgaluinb[17] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_nor02x1 \ALUSHT/ALU/U450  ( .ZN(\ALUSHT/ALU/pkaddina[1] ), .A(
        \ALUSHT/ALU/n1852 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_invx05 \ALUSHT/ALU/U589  ( .ZN(\ALUSHT/ALU/n1840 ), .A(\pgaluina[13] )
         );
    snl_xor2x0 \ALUSHT/ALU/U822  ( .Z(\ALUSHT/ALU/n2290 ), .A(
        \ALUSHT/ALU/intb[25] ), .B(\ALUSHT/ALU/intb[23] ) );
    snl_oai222x0 \ALUSHT/ALU/U477  ( .ZN(\ALUSHT/ALU/pkincin[6] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1894 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1847 ), .E(\ALUSHT/ALU/n1895 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nand04x0 \ALUSHT/ALU/U747  ( .ZN(\ALUSHT/ALU/n2257 ), .A(
        \ALUSHT/ALU/intb[23] ), .B(\ALUSHT/ALU/intb[24] ), .C(
        \ALUSHT/ALU/intb[25] ), .D(\ALUSHT/ALU/intb[26] ) );
    snl_ao022x1 \ALUSHT/ALU/U760  ( .Z(\ALUSHT/ALU/n2259 ), .A(
        \ALUSHT/ALU/pkdecout[8] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[8] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_ao022x1 \ALUSHT/ALU/U805  ( .Z(\ALUSHT/ALU/n2282 ), .A(
        \ALUSHT/ALU/pkdecout[16] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[16] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_muxi21x1 \ALUSHT/ALU/U995  ( .ZN(\ALUSHT/ALU/n1948 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1829 ) );
    snl_invx05 \ALUSHT/ALU/U577  ( .ZN(\ALUSHT/ALU/n1898 ), .A(\pgaluinb[4] )
         );
    snl_invx05 \ALUSHT/ALU/U895  ( .ZN(\ALUSHT/ALU/intb[21] ), .A(
        \ALUSHT/ALU/n1830 ) );
    snl_invx05 \ALUSHT/ALU/U905  ( .ZN(\ALUSHT/ALU/intb[18] ), .A(
        \ALUSHT/ALU/n1833 ) );
    snl_muxi21x1 \ALUSHT/ALU/U939  ( .ZN(\ALUSHT/ALU/n2162 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1894 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1025  ( .ZN(\ALUSHT/ALU/n1978 ), .A(
        \ALUSHT/ALU/n2236 ), .B(\ALUSHT/ALU/n2235 ), .S(\ALUSHT/ALU/n1839 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1002  ( .ZN(\ALUSHT/ALU/n1954 ), .A(
        \ALUSHT/ALU/n2210 ), .B(\ALUSHT/ALU/n2211 ), .S(\ALUSHT/ALU/inta[20] )
         );
    snl_nand13x2 \ALUSHT/ALU/U374  ( .ZN(\ALUSHT/ALU/n2103 ), .A(
        \ALUSHT/ALU/pkaddcin ), .B(\ALUSHT/ALU/n2119 ), .C(\ALUSHT/ALU/n1818 )
         );
    snl_nand02x2 \ALUSHT/ALU/U383  ( .ZN(\ALUSHT/ALU/n1857 ), .A(
        \ALUSHT/ALU/n2077 ), .B(\ALUSHT/ALU/n2078 ) );
    snl_nor02x1 \ALUSHT/ALU/U425  ( .ZN(\ALUSHT/ALU/pkaddina[27] ), .A(
        \ALUSHT/ALU/n1807 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U550  ( .ZN(\ALUSHT/ALU/n2054 ), .A(
        \ALUSHT/ALU/n2055 ), .B(\ALUSHT/ALU/n2056 ) );
    snl_nand03x0 \ALUSHT/ALU/U647  ( .ZN(\ALUSHT/ALU/n2175 ), .A(
        \ALUSHT/ALU/n2174 ), .B(\ALUSHT/ALU/n2152 ), .C(\ALUSHT/ALU/n2176 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1019  ( .ZN(\ALUSHT/ALU/n2227 ), .A(
        \ALUSHT/ALU/n2145 ), .B(\ALUSHT/ALU/n2143 ), .S(\ALUSHT/ALU/intb[16] )
         );
    snl_oai012x1 \ALUSHT/ALU/U660  ( .ZN(\ALUSHT/ALU/n2195 ), .A(
        \ALUSHT/ALU/intb[25] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_nand02x1 \ALUSHT/ALU/U922  ( .ZN(\ALUSHT/ALU/n1975 ), .A(
        \ALUSHT/ALU/pkaddsum[15] ), .B(\ALUSHT/ALU/n2103 ) );
    snl_mux21x1 \ALUSHT/ALU/U685  ( .Z(\ALUSHT/ALU/n2232 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2233 ), .S(\ALUSHT/ALU/n2091 ) );
    snl_nand12x1 \ALUSHT/ALU/U839  ( .ZN(\ALUSHT/ALU/n2101 ), .A(
        \ALUSHT/ALU/n2093 ), .B(\ALUSHT/ALU/n2078 ) );
    snl_muxi21x1 \ALUSHT/ALU/U715  ( .ZN(\ALUSHT/ALU/pkaddinb[25] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1826 ) );
    snl_nor02x1 \ALUSHT/ALU/U857  ( .ZN(\ALUSHT/ALU/n1901 ), .A(
        \ALUSHT/ALU/n1900 ), .B(\pgaluina[3] ) );
    snl_invx05 \ALUSHT/ALU/U870  ( .ZN(\ALUSHT/ALU/n2061 ), .A(
        \ALUSHT/ALU/n1861 ) );
    snl_aoi012x1 \ALUSHT/ALU/U391  ( .ZN(\ALUSHT/ALU/n1805 ), .A(
        \pgaluina[29] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U402  ( .ZN(\ALUSHT/ALU/n1816 ), .A(
        \pgaluina[18] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_nor02x1 \ALUSHT/ALU/U437  ( .ZN(\ALUSHT/ALU/pkaddina[14] ), .A(
        \ALUSHT/ALU/n1839 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U489  ( .ZN(\ALUSHT/ALU/pkdecin[25] ), .A(
        \ALUSHT/ALU/n1809 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_invx05 \ALUSHT/ALU/U592  ( .ZN(\ALUSHT/ALU/n1882 ), .A(\pgaluinb[12] )
         );
    snl_nor04x0 \ALUSHT/ALU/U732  ( .ZN(\ALUSHT/ALU/n2064 ), .A(
        \ALUSHT/ALU/n1864 ), .B(\ALUSHT/ALU/n1865 ), .C(\ALUSHT/ALU/n1866 ), 
        .D(\ALUSHT/ALU/n1867 ) );
    snl_xnor2x0 \ALUSHT/ALU/U1050  ( .ZN(\ALUSHT/ALU/n2294 ), .A(
        \ALUSHT/ALU/n1882 ), .B(\ALUSHT/ALU/n1880 ) );
    snl_nand04x0 \ALUSHT/ALU/U519  ( .ZN(\ALUSHT/pkaluout[26] ), .A(
        \ALUSHT/ALU/n1930 ), .B(\ALUSHT/ALU/n1931 ), .C(\ALUSHT/ALU/n1932 ), 
        .D(\ALUSHT/ALU/n1933 ) );
    snl_and08x1 \ALUSHT/ALU/U629  ( .Z(\ALUSHT/ALU/n2135 ), .A(\pgaluina[10] ), 
        .B(\pgaluina[11] ), .C(\pgaluina[0] ), .D(\ALUSHT/ALU/n2136 ), .E(
        \ALUSHT/ALU/n2137 ), .F(\pgaluina[9] ), .G(\ALUSHT/ALU/n2138 ), .H(
        \ALUSHT/ALU/n2139 ) );
    snl_oai012x1 \ALUSHT/ALU/U697  ( .ZN(\ALUSHT/ALU/n2250 ), .A(\pgaluinb[0] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U707  ( .ZN(\ALUSHT/ALU/pkaddinb[3] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[3] ) );
    snl_muxi21x1 \ALUSHT/ALU/U979  ( .ZN(\ALUSHT/ALU/n1932 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1825 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1042  ( .ZN(\ALUSHT/ALU/n2035 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1907 ) );
    snl_invx05 \ALUSHT/ALU/U580  ( .ZN(\ALUSHT/ALU/n1876 ), .A(\pgaluina[15] )
         );
    snl_nor02x1 \ALUSHT/ALU/U845  ( .ZN(\ALUSHT/ALU/n1804 ), .A(
        \ALUSHT/ALU/n1876 ), .B(\ALUSHT/ALU/n1803 ) );
    snl_aoi012x1 \ALUSHT/ALU/U410  ( .ZN(\ALUSHT/ALU/n1825 ), .A(
        \pgaluinb[26] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_oai222x0 \ALUSHT/ALU/U459  ( .ZN(\ALUSHT/ALU/pkincin[24] ), .A(
        \ALUSHT/ALU/n1827 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1810 ), .E(\ALUSHT/ALU/n1866 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_muxi21x1 \ALUSHT/ALU/U720  ( .ZN(\ALUSHT/ALU/pkaddinb[20] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1831 ) );
    snl_invx05 \ALUSHT/ALU/U862  ( .ZN(\ALUSHT/ALU/inta[30] ), .A(
        \ALUSHT/ALU/n1802 ) );
    snl_aoi112x0 \ALUSHT/ALU/U769  ( .ZN(\ALUSHT/ALU/n2021 ), .A(
        \ALUSHT/ALU/pkaddsum[4] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2263 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U442  ( .ZN(\ALUSHT/ALU/pkaddina[9] ), .A(
        \ALUSHT/ALU/n1844 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nand04x0 \ALUSHT/ALU/U542  ( .ZN(\ALUSHT/pkaluout[3] ), .A(
        \ALUSHT/ALU/n2022 ), .B(\ALUSHT/ALU/n2023 ), .C(\ALUSHT/ALU/n2024 ), 
        .D(\ALUSHT/ALU/n2025 ) );
    snl_invx05 \ALUSHT/ALU/U565  ( .ZN(\ALUSHT/ALU/n1888 ), .A(\pgaluinb[9] )
         );
    snl_nand02x1 \ALUSHT/ALU/U655  ( .ZN(\ALUSHT/ALU/n2187 ), .A(
        \ALUSHT/ALU/n2188 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nor02x1 \ALUSHT/ALU/U887  ( .ZN(\ALUSHT/ALU/n1866 ), .A(
        \ALUSHT/ALU/n1827 ), .B(\ALUSHT/ALU/inta[24] ) );
    snl_nor02x1 \ALUSHT/ALU/U917  ( .ZN(\ALUSHT/ALU/n1885 ), .A(
        \ALUSHT/ALU/n1884 ), .B(\pgaluina[11] ) );
    snl_oai012x1 \ALUSHT/ALU/U672  ( .ZN(\ALUSHT/ALU/n2213 ), .A(\pgaluinb[1] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_invx05 \ALUSHT/ALU/U559  ( .ZN(\ALUSHT/ALU/n2044 ), .A(\poalufnc[4] )
         );
    snl_muxi21x1 \ALUSHT/ALU/U930  ( .ZN(\ALUSHT/ALU/n1998 ), .A(
        \ALUSHT/ALU/n2147 ), .B(\ALUSHT/ALU/n2149 ), .S(\pgaluina[9] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1037  ( .ZN(\ALUSHT/ALU/n1992 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[11] ) );
    snl_nand02x1 \ALUSHT/ALU/U669  ( .ZN(\ALUSHT/ALU/n2208 ), .A(
        \ALUSHT/ALU/n2209 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1010  ( .ZN(\ALUSHT/ALU/n1960 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1832 ) );
    snl_oai222x0 \ALUSHT/ALU/U465  ( .ZN(\ALUSHT/ALU/pkincin[18] ), .A(
        \ALUSHT/ALU/n1833 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1816 ), .E(\ALUSHT/ALU/n1872 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nor02x1 \ALUSHT/ALU/U755  ( .ZN(\ALUSHT/ALU/n2138 ), .A(
        \ALUSHT/ALU/n1845 ), .B(\ALUSHT/ALU/n1846 ) );
    snl_ao022x1 \ALUSHT/ALU/U772  ( .Z(\ALUSHT/ALU/n2265 ), .A(
        \ALUSHT/ALU/pkdecout[31] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[31] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_invx05 \ALUSHT/ALU/U830  ( .ZN(\ALUSHT/ALU/n2084 ), .A(
        \ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U480  ( .ZN(\ALUSHT/ALU/pkincin[3] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1900 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1850 ), .E(\ALUSHT/ALU/n1901 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_and02x1 \ALUSHT/ALU/U510  ( .Z(\ALUSHT/ALU/pkdecin[3] ), .A(
        \pgaluina[3] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_muxi21x1 \ALUSHT/ALU/U620  ( .ZN(\ALUSHT/ALU/n2118 ), .A(
        \ALUSHT/ALU/n2058 ), .B(exetype1), .S(\ALUSHT/ALU/n1877 ) );
    snl_ao022x1 \ALUSHT/ALU/U817  ( .Z(\ALUSHT/ALU/n2287 ), .A(
        \ALUSHT/ALU/pkdecout[10] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[10] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_invx05 \ALUSHT/ALU/U879  ( .ZN(\ALUSHT/ALU/inta[26] ), .A(
        \ALUSHT/ALU/n1808 ) );
    snl_muxi21x1 \ALUSHT/ALU/U987  ( .ZN(\ALUSHT/ALU/n1940 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1827 ) );
    snl_nand04x0 \ALUSHT/ALU/U537  ( .ZN(\ALUSHT/pkaluout[8] ), .A(
        \ALUSHT/ALU/n2002 ), .B(\ALUSHT/ALU/n2003 ), .C(\ALUSHT/ALU/n2004 ), 
        .D(\ALUSHT/ALU/n2005 ) );
    snl_muxi21x1 \ALUSHT/ALU/U962  ( .ZN(\ALUSHT/ALU/n2027 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1903 ) );
    snl_nand02x1 \ALUSHT/ALU/U607  ( .ZN(\ALUSHT/ALU/n2093 ), .A(
        \ALUSHT/ALU/n2092 ), .B(\poalufnc[2] ) );
    snl_ao022x1 \ALUSHT/ALU/U797  ( .Z(\ALUSHT/ALU/n2278 ), .A(
        \ALUSHT/ALU/pkdecout[1] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[1] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_muxi21x1 \ALUSHT/ALU/U945  ( .ZN(\ALUSHT/ALU/n2016 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[5] ) );
    snl_muxi21x1 \ALUSHT/ALU/U368  ( .ZN(\ALUSHT/ALU/n2006 ), .A(
        \ALUSHT/ALU/n2157 ), .B(\ALUSHT/ALU/n2158 ), .S(\pgaluina[7] ) );
    snl_nor02x1 \ALUSHT/ALU/U487  ( .ZN(\ALUSHT/ALU/pkdecin[27] ), .A(
        \ALUSHT/ALU/n1807 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_nand14x0 \ALUSHT/ALU/U530  ( .ZN(\ALUSHT/pkaluout[15] ), .A(
        \ALUSHT/ALU/n1974 ), .B(\ALUSHT/ALU/n1975 ), .C(\ALUSHT/ALU/n1976 ), 
        .D(\ALUSHT/ALU/n1977 ) );
    snl_aoi012x1 \ALUSHT/ALU/U600  ( .ZN(\ALUSHT/ALU/pkcmpina[31] ), .A(
        \pgaluina[31] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U859  ( .ZN(\ALUSHT/ALU/pkcmpinb[31] ), .A(
        \pgaluinb[31] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_aoi112x0 \ALUSHT/ALU/U790  ( .ZN(\ALUSHT/ALU/n1945 ), .A(
        \ALUSHT/ALU/pkaddsum[23] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2274 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U942  ( .ZN(\ALUSHT/ALU/n2012 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[6] ) );
    snl_muxi21x1 \ALUSHT/ALU/U965  ( .ZN(\ALUSHT/ALU/n1919 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1861 ) );
    snl_nand04x0 \ALUSHT/ALU/U517  ( .ZN(\ALUSHT/pkaluout[28] ), .A(
        \ALUSHT/ALU/n1922 ), .B(\ALUSHT/ALU/n1923 ), .C(\ALUSHT/ALU/n1924 ), 
        .D(\ALUSHT/ALU/n1925 ) );
    snl_invx05 \ALUSHT/ALU/U579  ( .ZN(\ALUSHT/ALU/n1900 ), .A(\pgaluinb[3] )
         );
    snl_or08x1 \ALUSHT/ALU/U627  ( .Z(\ALUSHT/ALU/n2130 ), .A(
        \ALUSHT/ALU/inta[30] ), .B(\ALUSHT/ALU/inta[29] ), .C(
        \ALUSHT/ALU/inta[28] ), .D(\ALUSHT/ALU/inta[27] ), .E(
        \ALUSHT/ALU/inta[26] ), .F(\ALUSHT/ALU/n2131 ), .G(\ALUSHT/ALU/n2132 ), 
        .H(\ALUSHT/ALU/n2133 ) );
    snl_nand03x2 \ALUSHT/ALU/U373  ( .ZN(\ALUSHT/ALU/n1836 ), .A(
        \ALUSHT/ALU/n2073 ), .B(\ALUSHT/ALU/n2045 ), .C(\poalufnc[4] ) );
    snl_nor02x1 \ALUSHT/ALU/U445  ( .ZN(\ALUSHT/ALU/pkaddina[6] ), .A(
        \ALUSHT/ALU/n1847 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U462  ( .ZN(\ALUSHT/ALU/pkincin[21] ), .A(
        \ALUSHT/ALU/n1830 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1813 ), .E(\ALUSHT/ALU/n1869 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nand02x1 \ALUSHT/ALU/U649  ( .ZN(\ALUSHT/ALU/n2178 ), .A(
        \ALUSHT/ALU/n2179 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1017  ( .ZN(\ALUSHT/ALU/n1966 ), .A(
        \ALUSHT/ALU/n2222 ), .B(\ALUSHT/ALU/n2223 ), .S(\ALUSHT/ALU/inta[17] )
         );
    snl_aoi112x0 \ALUSHT/ALU/U810  ( .ZN(\ALUSHT/ALU/n1981 ), .A(
        \ALUSHT/ALU/pkaddsum[14] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2283 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U980  ( .ZN(\ALUSHT/ALU/n2197 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1826 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1030  ( .ZN(\ALUSHT/ALU/n1984 ), .A(
        \ALUSHT/ALU/n2151 ), .B(\ALUSHT/ALU/n2153 ), .S(\pgaluinb[13] ) );
    snl_nor04x0 \ALUSHT/ALU/U752  ( .ZN(\ALUSHT/ALU/n2128 ), .A(
        \ALUSHT/ALU/n1810 ), .B(\ALUSHT/ALU/n1808 ), .C(\ALUSHT/ALU/n1809 ), 
        .D(\ALUSHT/ALU/n1811 ) );
    snl_aoi112x0 \ALUSHT/ALU/U775  ( .ZN(\ALUSHT/ALU/n1917 ), .A(
        \ALUSHT/ALU/pkaddsum[30] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2266 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nand12x1 \ALUSHT/ALU/U837  ( .ZN(\ALUSHT/ALU/n2144 ), .A(
        \ALUSHT/ALU/n2046 ), .B(\ALUSHT/ALU/n2083 ) );
    snl_oai222x0 \ALUSHT/ALU/U479  ( .ZN(\ALUSHT/ALU/pkincin[4] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1898 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1849 ), .E(\ALUSHT/ALU/n1899 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_and05x1 \ALUSHT/ALU/U749  ( .Z(\ALUSHT/ALU/n2051 ), .A(
        \ALUSHT/ALU/intb[21] ), .B(\ALUSHT/ALU/intb[22] ), .C(
        \ALUSHT/ALU/intb[20] ), .D(\ALUSHT/ALU/intb[18] ), .E(
        \ALUSHT/ALU/intb[19] ) );
    snl_nand04x0 \ALUSHT/ALU/U545  ( .ZN(\ALUSHT/pkaluout[0] ), .A(
        \ALUSHT/ALU/n2034 ), .B(\ALUSHT/ALU/n2035 ), .C(\ALUSHT/ALU/n2036 ), 
        .D(\ALUSHT/ALU/n2037 ) );
    snl_muxi21x1 \ALUSHT/ALU/U937  ( .ZN(\ALUSHT/ALU/n2007 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1893 ) );
    snl_and02x1 \ALUSHT/ALU/U562  ( .Z(\ALUSHT/ALU/n2077 ), .A(\poalufnc[4] ), 
        .B(\ALUSHT/ALU/n2074 ) );
    snl_oai012x1 \ALUSHT/ALU/U652  ( .ZN(\ALUSHT/ALU/n2183 ), .A(
        \ALUSHT/ALU/intb[29] ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 )
         );
    snl_nand02x1 \ALUSHT/ALU/U675  ( .ZN(\ALUSHT/ALU/n2217 ), .A(
        \ALUSHT/ALU/n2218 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_invx05 \ALUSHT/ALU/U880  ( .ZN(\ALUSHT/ALU/intb[26] ), .A(
        \ALUSHT/ALU/n1825 ) );
    snl_invx05 \ALUSHT/ALU/U910  ( .ZN(\ALUSHT/ALU/n1838 ), .A(
        \ALUSHT/ALU/inta[16] ) );
    snl_nand02x2 \ALUSHT/ALU/U384  ( .ZN(\ALUSHT/ALU/n1860 ), .A(
        \ALUSHT/ALU/n2080 ), .B(\ALUSHT/ALU/n2077 ) );
    snl_aoi012x1 \ALUSHT/ALU/U396  ( .ZN(\ALUSHT/ALU/n1810 ), .A(
        \pgaluina[24] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1804 ) );
    snl_aoi012x1 \ALUSHT/ALU/U417  ( .ZN(\ALUSHT/ALU/n1832 ), .A(
        \pgaluinb[19] ), .B(\ALUSHT/ALU/n1803 ), .C(\ALUSHT/ALU/n1821 ) );
    snl_muxi21x1 \ALUSHT/ALU/U727  ( .ZN(\ALUSHT/ALU/pkaddinb[13] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\pgaluinb[13] ) );
    snl_muxi21x1 \ALUSHT/ALU/U959  ( .ZN(\ALUSHT/ALU/n1914 ), .A(
        \ALUSHT/ALU/n2177 ), .B(\ALUSHT/ALU/n2178 ), .S(\ALUSHT/ALU/inta[30] )
         );
    snl_xor2x0 \ALUSHT/ALU/U1045  ( .Z(\ALUSHT/ALU/n2108 ), .A(
        \ALUSHT/ALU/intb[29] ), .B(\ALUSHT/ALU/n1823 ) );
    snl_invx05 \ALUSHT/ALU/U865  ( .ZN(\ALUSHT/ALU/n2059 ), .A(
        \ALUSHT/ALU/n1859 ) );
    snl_oai012x1 \ALUSHT/ALU/U405  ( .ZN(\ALUSHT/ALU/pkaddcin ), .A(
        \ALUSHT/ALU/n1817 ), .B(\ALUSHT/ALU/n1818 ), .C(\ALUSHT/ALU/n1819 ) );
    snl_nor02x1 \ALUSHT/ALU/U430  ( .ZN(\ALUSHT/ALU/pkaddina[22] ), .A(
        \ALUSHT/ALU/n1812 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_invx05 \ALUSHT/ALU/U587  ( .ZN(\ALUSHT/ALU/n1839 ), .A(\pgaluina[14] )
         );
    snl_invx05 \ALUSHT/ALU/U842  ( .ZN(\ALUSHT/ALU/n2053 ), .A(
        \ALUSHT/ALU/n2081 ) );
    snl_invx05 \ALUSHT/ALU/U595  ( .ZN(\ALUSHT/ALU/n1843 ), .A(\pgaluina[10] )
         );
    snl_nand02x1 \ALUSHT/ALU/U690  ( .ZN(\ALUSHT/ALU/n2239 ), .A(
        \ALUSHT/ALU/n2240 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U700  ( .ZN(\ALUSHT/ALU/n2043 ), .A(
        \ALUSHT/ALU/n2254 ), .B(\ALUSHT/ALU/n2067 ), .S(\poalufnc[2] ) );
    snl_or05x1 \ALUSHT/ALU/U735  ( .Z(\ALUSHT/ALU/n2039 ), .A(
        \ALUSHT/ALU/n1889 ), .B(\ALUSHT/ALU/n1891 ), .C(\ALUSHT/ALU/n1893 ), 
        .D(\ALUSHT/ALU/n1895 ), .E(\ALUSHT/ALU/n1897 ) );
    snl_nor02x1 \ALUSHT/ALU/U422  ( .ZN(\ALUSHT/ALU/pkaddina[30] ), .A(
        \ALUSHT/ALU/n1802 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_nor02x1 \ALUSHT/ALU/U877  ( .ZN(\ALUSHT/ALU/n1863 ), .A(
        \ALUSHT/ALU/inta[27] ), .B(\ALUSHT/ALU/n1824 ) );
    snl_nor02x1 \ALUSHT/ALU/U439  ( .ZN(\ALUSHT/ALU/pkaddina[12] ), .A(
        \ALUSHT/ALU/n1841 ), .B(\ALUSHT/ALU/n1836 ) );
    snl_oai222x0 \ALUSHT/ALU/U457  ( .ZN(\ALUSHT/ALU/pkincin[26] ), .A(
        \ALUSHT/ALU/n1825 ), .B(\ALUSHT/ALU/n1857 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1808 ), .E(\ALUSHT/ALU/n1864 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_oai222x0 \ALUSHT/ALU/U470  ( .ZN(\ALUSHT/ALU/pkincin[13] ), .A(
        \ALUSHT/ALU/n1857 ), .B(\ALUSHT/ALU/n1880 ), .C(\ALUSHT/ALU/n1858 ), 
        .D(\ALUSHT/ALU/n1840 ), .E(\ALUSHT/ALU/n1881 ), .F(\ALUSHT/ALU/n1860 )
         );
    snl_nand04x0 \ALUSHT/ALU/U539  ( .ZN(\ALUSHT/pkaluout[6] ), .A(
        \ALUSHT/ALU/n2010 ), .B(\ALUSHT/ALU/n2011 ), .C(\ALUSHT/ALU/n2012 ), 
        .D(\ALUSHT/ALU/n2013 ) );
    snl_muxi21x1 \ALUSHT/ALU/U682  ( .ZN(\ALUSHT/ALU/n2056 ), .A(
        \ALUSHT/ALU/n2148 ), .B(\ALUSHT/ALU/n2228 ), .S(\pgaluina[15] ) );
    snl_muxi21x1 \ALUSHT/ALU/U712  ( .ZN(\ALUSHT/ALU/pkaddinb[28] ), .A(
        \ALUSHT/ALU/n2069 ), .B(\ALUSHT/ALU/n1818 ), .S(\ALUSHT/ALU/intb[28] )
         );
    snl_invx05 \ALUSHT/ALU/U850  ( .ZN(\ALUSHT/ALU/n2078 ), .A(
        \ALUSHT/ALU/n2075 ) );
    snl_invx05 \ALUSHT/ALU/U557  ( .ZN(\ALUSHT/ALU/n2073 ), .A(\poalufnc[2] )
         );
    snl_nor03x0 \ALUSHT/ALU/U609  ( .ZN(\ALUSHT/ALU/n2096 ), .A(\poalufnc[3] ), 
        .B(\poalufnc[4] ), .C(\poalufnc[2] ) );
    snl_ao022x1 \ALUSHT/ALU/U799  ( .Z(\ALUSHT/ALU/n2279 ), .A(
        \ALUSHT/ALU/pkdecout[19] ), .B(\ALUSHT/ALU/n2105 ), .C(
        \ALUSHT/ALU/pkincout[19] ), .D(\ALUSHT/ALU/n2104 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1039  ( .ZN(\ALUSHT/ALU/n1995 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1887 ) );
    snl_invx05 \ALUSHT/ALU/U570  ( .ZN(\ALUSHT/ALU/n1846 ), .A(\pgaluina[7] )
         );
    snl_nand02x1 \ALUSHT/ALU/U640  ( .ZN(\ALUSHT/ALU/n2164 ), .A(
        \ALUSHT/ALU/n2165 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_nand02x1 \ALUSHT/ALU/U667  ( .ZN(\ALUSHT/ALU/n2205 ), .A(
        \ALUSHT/ALU/n2206 ), .B(\ALUSHT/ALU/n2100 ) );
    snl_muxi21x1 \ALUSHT/ALU/U925  ( .ZN(\ALUSHT/ALU/n2122 ), .A(
        \ALUSHT/ALU/n2120 ), .B(\ALUSHT/ALU/n2121 ), .S(
        \ALUSHT/ALU/pkaddina[15] ) );
    snl_ao022x1 \ALUSHT/ALU/U819  ( .Z(\ALUSHT/ALU/n2288 ), .A(
        \ALUSHT/ALU/pkdecout[0] ), .B(\ALUSHT/ALU/n1909 ), .C(
        \ALUSHT/ALU/pkincout[0] ), .D(\ALUSHT/ALU/n1855 ) );
    snl_invx05 \ALUSHT/ALU/U892  ( .ZN(\ALUSHT/ALU/intb[22] ), .A(
        \ALUSHT/ALU/n1829 ) );
    snl_invx05 \ALUSHT/ALU/U902  ( .ZN(\ALUSHT/ALU/intb[19] ), .A(
        \ALUSHT/ALU/n1832 ) );
    snl_muxi21x1 \ALUSHT/ALU/U989  ( .ZN(\ALUSHT/ALU/n1943 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1867 ) );
    snl_nand04x0 \ALUSHT/ALU/U740  ( .ZN(\ALUSHT/ALU/n2133 ), .A(
        \ALUSHT/ALU/pkdecin[31] ), .B(\ALUSHT/ALU/n1876 ), .C(
        \ALUSHT/ALU/n1838 ), .D(\ALUSHT/ALU/n1837 ) );
    snl_aoi112x0 \ALUSHT/ALU/U802  ( .ZN(\ALUSHT/ALU/n1965 ), .A(
        \ALUSHT/ALU/pkaddsum[18] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2280 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_muxi21x1 \ALUSHT/ALU/U992  ( .ZN(\ALUSHT/ALU/n2206 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1829 ) );
    snl_aoi112x0 \ALUSHT/ALU/U767  ( .ZN(\ALUSHT/ALU/n2017 ), .A(
        \ALUSHT/ALU/pkaddsum[5] ), .B(\ALUSHT/ALU/n2103 ), .C(
        \ALUSHT/ALU/n2262 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_nor02x1 \ALUSHT/ALU/U495  ( .ZN(\ALUSHT/ALU/pkdecin[19] ), .A(
        \ALUSHT/ALU/n1815 ), .B(\ALUSHT/ALU/n1908 ) );
    snl_and02x1 \ALUSHT/ALU/U505  ( .Z(\ALUSHT/ALU/pkdecin[8] ), .A(
        \pgaluina[8] ), .B(\ALUSHT/ALU/n1909 ) );
    snl_nand04x0 \ALUSHT/ALU/U522  ( .ZN(\ALUSHT/pkaluout[23] ), .A(
        \ALUSHT/ALU/n1942 ), .B(\ALUSHT/ALU/n1943 ), .C(\ALUSHT/ALU/n1944 ), 
        .D(\ALUSHT/ALU/n1945 ) );
    snl_oa012x1 \ALUSHT/ALU/U612  ( .Z(\ALUSHT/ALU/n2100 ), .A(
        \ALUSHT/ALU/n2079 ), .B(\ALUSHT/ALU/n2093 ), .C(\ALUSHT/ALU/n2101 ) );
    snl_aoi112x0 \ALUSHT/ALU/U782  ( .ZN(\ALUSHT/ALU/n1929 ), .A(
        \ALUSHT/ALU/pkaddsum[27] ), .B(\ALUSHT/ALU/n2102 ), .C(
        \ALUSHT/ALU/n2270 ), .D(\ALUSHT/ALU/n1974 ) );
    snl_xor3x1 \ALUSHT/ALU/U825  ( .Z(\ALUSHT/ALU/n2114 ), .A(
        \ALUSHT/ALU/n2109 ), .B(\ALUSHT/ALU/intb[16] ), .C(\ALUSHT/ALU/n2294 )
         );
    snl_invx05 \ALUSHT/ALU/U889  ( .ZN(\ALUSHT/ALU/intb[23] ), .A(
        \ALUSHT/ALU/n1828 ) );
    snl_nor02x1 \ALUSHT/ALU/U919  ( .ZN(\ALUSHT/ALU/n1907 ), .A(
        \ALUSHT/ALU/n1906 ), .B(\pgaluina[0] ) );
    snl_muxi21x1 \ALUSHT/ALU/U1005  ( .ZN(\ALUSHT/ALU/n2031 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1905 ) );
    snl_muxi21x1 \ALUSHT/ALU/U1022  ( .ZN(\ALUSHT/ALU/n1972 ), .A(
        \ALUSHT/ALU/n2153 ), .B(\ALUSHT/ALU/n2151 ), .S(\ALUSHT/ALU/n1835 ) );
    snl_muxi21x1 \ALUSHT/ALU/U950  ( .ZN(\ALUSHT/ALU/n2171 ), .A(
        \ALUSHT/ALU/n2143 ), .B(\ALUSHT/ALU/n2145 ), .S(\ALUSHT/ALU/n1900 ) );
    snl_oai012x1 \ALUSHT/ALU/U635  ( .ZN(\ALUSHT/ALU/n2157 ), .A(\pgaluinb[7] 
        ), .B(\ALUSHT/ALU/n2148 ), .C(\ALUSHT/ALU/n2097 ) );
    snl_muxi21x1 \ALUSHT/ALU/U977  ( .ZN(\ALUSHT/ALU/n1931 ), .A(
        \ALUSHT/ALU/n2296 ), .B(\ALUSHT/ALU/n2095 ), .S(\ALUSHT/ALU/n1864 ) );
    snl_muxi21x1 \ALUSHT/ALU/U699  ( .ZN(\ALUSHT/ALU/n2253 ), .A(
        \ALUSHT/ALU/pkgtflg ), .B(\ALUSHT/ALU/n2057 ), .S(\poalufnc[1] ) );
    snl_muxi21x1 \ALUSHT/ALU/U709  ( .ZN(\ALUSHT/ALU/pkaddinb[30] ), .A(
        \ALUSHT/ALU/n1818 ), .B(\ALUSHT/ALU/n2069 ), .S(\ALUSHT/ALU/n1820 ) );
    snl_aoi022x1 \ALUSHT/SHT/U274  ( .ZN(\ALUSHT/SHT/n2387 ), .A(
        \pgaluina[31] ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2389 ), .D(
        \ALUSHT/SHT/n2390 ) );
    snl_oa2222x1 \ALUSHT/SHT/U275  ( .Z(\ALUSHT/SHT/n2396 ), .A(
        \ALUSHT/SHT/n2397 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2398 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2400 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2401 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_oa2222x1 \ALUSHT/SHT/U276  ( .Z(\ALUSHT/SHT/n2545 ), .A(
        \ALUSHT/SHT/n2926 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2927 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2929 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2928 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_oa2222x1 \ALUSHT/SHT/U278  ( .Z(\ALUSHT/SHT/n2588 ), .A(
        \ALUSHT/SHT/n2922 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2923 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2925 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2924 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U286  ( .ZN(\ALUSHT/SHT/n2385 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[2] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[3] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[4] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[1] ) );
    snl_aoi122x0 \ALUSHT/SHT/U294  ( .ZN(\ALUSHT/SHT/n2966 ), .A(
        \pgaluina[14] ), .B(\ALUSHT/SHT/n2915 ), .C(\ALUSHT/SHT/n2965 ), .D(
        \phshtd[4] ), .E(\ALUSHT/SHT/n2492 ) );
    snl_aoi022x1 \ALUSHT/SHT/U304  ( .ZN(\ALUSHT/SHT/n2551 ), .A(
        \ALUSHT/SHT/n2541 ), .B(\pgaluina[0] ), .C(\ALUSHT/SHT/n2506 ), .D(
        \pgaluina[1] ) );
    snl_aoi122x0 \ALUSHT/SHT/U338  ( .ZN(\ALUSHT/SHT/n2349 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[15] ), .C(\pgaluina[23] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi022x4 \ALUSHT/SHT/U394  ( .ZN(\ALUSHT/SHT/n2647 ), .A(
        \pgaluina[12] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[11] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi2222x2 \ALUSHT/SHT/U415  ( .ZN(\ALUSHT/SHT/n2328 ), .A(
        \ALUSHT/SHT/n2660 ), .B(\ALUSHT/SHT/n2893 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2894 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[4] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2895 ) );
    snl_aoi012x4 \ALUSHT/SHT/U432  ( .ZN(\ALUSHT/SHT/n2699 ), .A(
        \ALUSHT/SHT/n2694 ), .B(\ALUSHT/SHT/n2700 ), .C(\ALUSHT/SHT/n2696 ) );
    snl_ao012x1 \ALUSHT/SHT/U692  ( .Z(\ALUSHT/SHT/n2471 ), .A(\pgaluina[1] ), 
        .B(\ALUSHT/SHT/n2651 ), .C(\ALUSHT/SHT/n2492 ) );
    snl_aoi012x1 \ALUSHT/SHT/U840  ( .ZN(\ALUSHT/SHT/n2985 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[23] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_invx05 \ALUSHT/SHT/U702  ( .ZN(\ALUSHT/SHT/n2477 ), .A(
        \ALUSHT/SHT/n2374 ) );
    snl_nand02x1 \ALUSHT/SHT/U725  ( .ZN(\ALUSHT/SHT/n2912 ), .A(
        \ALUSHT/SHT/n2909 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_invx05 \ALUSHT/SHT/U529  ( .ZN(\ALUSHT/SHT/n2381 ), .A(exetype1) );
    snl_oai122x0 \ALUSHT/SHT/U585  ( .ZN(\ALUSHT/SHT/n2605 ), .A(
        \ALUSHT/SHT/n2577 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2576 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi022x1 \ALUSHT/SHT/U867  ( .ZN(\ALUSHT/SHT/n3007 ), .A(
        \pgaluina[28] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[27] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U356  ( .ZN(\ALUSHT/SHT/n2314 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2743 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2744 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[13] ), 
        .G(\ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2745 ) );
    snl_invx1 \ALUSHT/SHT/U371  ( .ZN(\ALUSHT/SHT/n2682 ), .A(
        \ALUSHT/SHT/n2619 ) );
    snl_nor02x1 \ALUSHT/SHT/U560  ( .ZN(\ALUSHT/SHT/n2542 ), .A(
        \ALUSHT/SHT/n2522 ), .B(\ALUSHT/SHT/n2499 ) );
    snl_and02x1 \ALUSHT/SHT/U619  ( .Z(\ALUSHT/SHT/n2643 ), .A(
        \ALUSHT/SHT/n2622 ), .B(\ALUSHT/SHT/n2381 ) );
    snl_oai122x0 \ALUSHT/SHT/U1047  ( .ZN(\ALUSHT/SHT/n2844 ), .A(
        \ALUSHT/SHT/n2566 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3044 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2842 ) );
    snl_or04x1 \ALUSHT/SHT/U650  ( .Z(\ALUSHT/SHT/n2704 ), .A(
        \ALUSHT/SHT/n2567 ), .B(\ALUSHT/SHT/n2563 ), .C(\ALUSHT/SHT/n2560 ), 
        .D(\ALUSHT/SHT/n2556 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U789  ( .ZN(\ALUSHT/SHT/n2937 ), .A(
        \ALUSHT/SHT/n2853 ), .B(\ALUSHT/SHT/n2298 ), .C(\ALUSHT/SHT/n2534 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1060  ( .ZN(\ALUSHT/SHT/n2865 ), .A(
        \ALUSHT/SHT/n3104 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3097 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3099 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3102 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai2222x0 \ALUSHT/SHT/U882  ( .ZN(\ALUSHT/SHT/n2729 ), .A(
        \ALUSHT/SHT/n2955 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n2958 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n3017 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n2950 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_aoi122x0 \ALUSHT/SHT/U912  ( .ZN(\ALUSHT/SHT/n3034 ), .A(
        \ALUSHT/SHT/n3033 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2881 ), 
        .D(\ALUSHT/SHT/n2298 ), .E(\ALUSHT/SHT/n2391 ) );
    snl_aoi222x1 \ALUSHT/SHT/U447  ( .ZN(\ALUSHT/SHT/n2817 ), .A(
        \ALUSHT/SHT/n2548 ), .B(\ALUSHT/SHT/n2790 ), .C(\ALUSHT/SHT/n2659 ), 
        .D(\ALUSHT/SHT/n2818 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2819 )
         );
    snl_invx05 \ALUSHT/SHT/U547  ( .ZN(\ALUSHT/SHT/n2414 ), .A(\pgaluina[3] )
         );
    snl_aoi012x1 \ALUSHT/SHT/U677  ( .ZN(\ALUSHT/SHT/n2773 ), .A(
        \ALUSHT/SHT/n2423 ), .B(\pgaluina[26] ), .C(\ALUSHT/SHT/n2419 ) );
    snl_oai2222x0 \ALUSHT/SHT/U935  ( .ZN(\ALUSHT/SHT/n2745 ), .A(
        \ALUSHT/SHT/n2691 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2996 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3001 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3028 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1029  ( .ZN(\ALUSHT/SHT/n2816 ), .A(
        \ALUSHT/SHT/n3091 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2678 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3066 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3086 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_invx05 \ALUSHT/SHT/U777  ( .ZN(\ALUSHT/SHT/n2552 ), .A(
        \ALUSHT/SHT/n2868 ) );
    snl_oai012x1 \ALUSHT/SHT/U809  ( .ZN(\ALUSHT/SHT/n2681 ), .A(
        \ALUSHT/SHT/n2518 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_ao022x1 \ALUSHT/SHT/U999  ( .Z(\ALUSHT/SHT/n2781 ), .A(
        \ALUSHT/SHT/n2445 ), .B(\pgaluina[31] ), .C(\ALUSHT/SHT/n2444 ), .D(
        \ALUSHT/SHT/n3076 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1085  ( .ZN(\ALUSHT/SHT/n2904 ), .A(
        \ALUSHT/SHT/n3093 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3094 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n3083 ), .F(\ALUSHT/SHT/n2642 ), 
        .G(\ALUSHT/SHT/n3082 ), .H(\ALUSHT/SHT/n2454 ) );
    snl_invx05 \ALUSHT/SHT/U1115  ( .ZN(\ALUSHT/SHT/n2970 ), .A(
        \ALUSHT/SHT/n2968 ) );
    snl_aoi222x2 \ALUSHT/SHT/U460  ( .ZN(\ALUSHT/SHT/n2876 ), .A(
        \ALUSHT/SHT/n2849 ), .B(\ALUSHT/SHT/n2835 ), .C(\ALUSHT/SHT/n2810 ), 
        .D(\ALUSHT/SHT/n2767 ), .E(\ALUSHT/SHT/n2662 ), .F(\ALUSHT/SHT/n2877 )
         );
    snl_aoi012x1 \ALUSHT/SHT/U835  ( .ZN(\ALUSHT/SHT/n2448 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[18] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_nand02x1 \ALUSHT/SHT/U485  ( .ZN(\ALUSHT/pkshtout[19] ), .A(
        \ALUSHT/SHT/n2341 ), .B(\ALUSHT/SHT/n2342 ) );
    snl_invx05 \ALUSHT/SHT/U750  ( .ZN(\ALUSHT/SHT/n2702 ), .A(
        \ALUSHT/SHT/n2398 ) );
    snl_oai012x1 \ALUSHT/SHT/U812  ( .ZN(\ALUSHT/SHT/n2431 ), .A(
        \ALUSHT/SHT/n2519 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_oa122x1 \ALUSHT/SHT/U982  ( .Z(\ALUSHT/SHT/n2676 ), .A(
        \ALUSHT/SHT/n3068 ), .B(\ALUSHT/SHT/n2627 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n3067 ), .E(\ALUSHT/SHT/n2773 ) );
    snl_invx05 \ALUSHT/SHT/U899  ( .ZN(\ALUSHT/SHT/n3028 ), .A(
        \ALUSHT/SHT/n3027 ) );
    snl_oai2222x0 \ALUSHT/SHT/U909  ( .ZN(\ALUSHT/SHT/n2881 ), .A(
        \ALUSHT/SHT/n3006 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3010 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3008 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3007 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_invx05 \ALUSHT/SHT/U1015  ( .ZN(\ALUSHT/SHT/n2464 ), .A(
        \ALUSHT/SHT/n2486 ) );
    snl_oai122x0 \ALUSHT/SHT/U1032  ( .ZN(\ALUSHT/SHT/n2820 ), .A(
        \ALUSHT/SHT/n2582 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3093 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2817 ) );
    snl_oai122x0 \ALUSHT/SHT/U515  ( .ZN(\ALUSHT/SHT/n2447 ), .A(
        \ALUSHT/SHT/n2382 ), .B(\ALUSHT/SHT/n2448 ), .C(\ALUSHT/SHT/n2413 ), 
        .D(\ALUSHT/SHT/n2449 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_oa2222x1 \ALUSHT/SHT/U323  ( .Z(\ALUSHT/SHT/n2574 ), .A(
        \ALUSHT/SHT/n2928 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2929 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2531 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2930 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_invx05 \ALUSHT/SHT/U532  ( .ZN(\ALUSHT/SHT/n2366 ), .A(\pgaluina[31] )
         );
    snl_nand02x1 \ALUSHT/SHT/U602  ( .ZN(\ALUSHT/SHT/n2627 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n2382 ) );
    snl_oa022x1 \ALUSHT/SHT/U625  ( .Z(\ALUSHT/SHT/n2573 ), .A(
        \ALUSHT/SHT/n2532 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2558 ), 
        .D(\ALUSHT/SHT/n2399 ) );
    snl_oai012x1 \ALUSHT/SHT/U967  ( .ZN(\ALUSHT/SHT/n2417 ), .A(
        \ALUSHT/SHT/n2512 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_aoi022x1 \ALUSHT/SHT/U792  ( .ZN(\ALUSHT/SHT/n2940 ), .A(
        \pgaluina[21] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[20] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi012x4 \ALUSHT/SHT/U429  ( .ZN(\ALUSHT/SHT/n2697 ), .A(
        \ALUSHT/SHT/n2694 ), .B(\ALUSHT/SHT/n2698 ), .C(\ALUSHT/SHT/n2696 ) );
    snl_aoi222x0 \ALUSHT/SHT/U689  ( .ZN(\ALUSHT/SHT/n2348 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2840 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2841 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2837 )
         );
    snl_oa122x1 \ALUSHT/SHT/U940  ( .Z(\ALUSHT/SHT/n3051 ), .A(
        \ALUSHT/SHT/n3003 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n2648 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2384 ) );
    snl_invx05 \ALUSHT/SHT/U719  ( .ZN(\ALUSHT/SHT/n2663 ), .A(
        \ALUSHT/SHT/n2501 ) );
    snl_aoi012x1 \ALUSHT/SHT/U507  ( .ZN(\ALUSHT/SHT/n2406 ), .A(
        \ALUSHT/SHT/n2404 ), .B(\ALUSHT/SHT/n2407 ), .C(\ALUSHT/SHT/n2394 ) );
    snl_oai012x1 \ALUSHT/SHT/U849  ( .ZN(\ALUSHT/SHT/n2995 ), .A(
        \ALUSHT/SHT/n2414 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_invx05 \ALUSHT/SHT/U975  ( .ZN(\ALUSHT/SHT/n3066 ), .A(
        \ALUSHT/SHT/n3065 ) );
    snl_oai223x0 \ALUSHT/SHT/U1069  ( .ZN(\ALUSHT/SHT/n2883 ), .A(
        \ALUSHT/SHT/n2504 ), .B(\phshtd[5] ), .C(\ALUSHT/SHT/n3075 ), .D(
        \ALUSHT/SHT/n3108 ), .E(\ALUSHT/SHT/n2629 ), .F(\ALUSHT/SHT/n3071 ), 
        .G(\ALUSHT/SHT/n2630 ) );
    snl_aoi022x1 \ALUSHT/SHT/U316  ( .ZN(\ALUSHT/SHT/n2674 ), .A(\pgaluina[6] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[5] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_ao1b1b2x0 \ALUSHT/SHT/U497  ( .Z(\ALUSHT/pkshtout[31] ), .A(
        \ALUSHT/SHT/n2365 ), .B(\ALUSHT/SHT/n2366 ), .C(\ALUSHT/SHT/n2368 ), 
        .D(\ALUSHT/SHT/n2367 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U331  ( .ZN(\ALUSHT/SHT/n3017 ), .A(
        \ALUSHT/SHT/n2685 ), .B(\ALUSHT/SHT/n2539 ), .C(\ALUSHT/SHT/n2946 ), 
        .D(\ALUSHT/SHT/n2404 ), .E(\ALUSHT/SHT/n2778 ), .F(\ALUSHT/SHT/n2390 ), 
        .G(\ALUSHT/SHT/n2945 ), .H(\ALUSHT/SHT/n2694 ) );
    snl_and02x1 \ALUSHT/SHT/U610  ( .Z(\ALUSHT/SHT/n2634 ), .A(
        \ALUSHT/SHT/n2633 ), .B(exetype1) );
    snl_nand03x0 \ALUSHT/SHT/U637  ( .ZN(\ALUSHT/SHT/n2379 ), .A(
        \ALUSHT/SHT/n2661 ), .B(\ALUSHT/SHT/n2504 ), .C(\ALUSHT/SHT/n2662 ) );
    snl_invx05 \ALUSHT/SHT/U780  ( .ZN(\ALUSHT/SHT/n2452 ), .A(
        \ALUSHT/SHT/n2494 ) );
    snl_invx05 \ALUSHT/SHT/U952  ( .ZN(\ALUSHT/SHT/n3052 ), .A(
        \ALUSHT/SHT/n2812 ) );
    snl_invx1 \ALUSHT/SHT/U378  ( .ZN(\ALUSHT/SHT/n2302 ), .A(
        \ALUSHT/SHT/n2661 ) );
    snl_aoi012x1 \ALUSHT/SHT/U520  ( .ZN(\ALUSHT/SHT/n2474 ), .A(
        \ALUSHT/SHT/n2390 ), .B(\ALUSHT/SHT/n2407 ), .C(\ALUSHT/SHT/n2475 ) );
    snl_oai223x0 \ALUSHT/SHT/U1007  ( .ZN(\ALUSHT/SHT/n2794 ), .A(
        \ALUSHT/SHT/n2392 ), .B(\ALUSHT/SHT/n3030 ), .C(\ALUSHT/SHT/n2502 ), 
        .D(\ALUSHT/SHT/n3080 ), .E(\ALUSHT/SHT/n2455 ), .F(\ALUSHT/SHT/n3079 ), 
        .G(\ALUSHT/SHT/n2451 ) );
    snl_oa222x1 \ALUSHT/SHT/U1020  ( .Z(\ALUSHT/SHT/n3086 ), .A(
        \ALUSHT/SHT/n2770 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2987 ), 
        .D(\ALUSHT/SHT/n2501 ), .E(\ALUSHT/SHT/n2769 ), .F(\ALUSHT/SHT/n2427 )
         );
    snl_aoi222x1 \ALUSHT/SHT/U455  ( .ZN(\ALUSHT/SHT/n2822 ), .A(
        \ALUSHT/SHT/n2548 ), .B(\ALUSHT/SHT/n2823 ), .C(\ALUSHT/SHT/n2659 ), 
        .D(\ALUSHT/SHT/n2824 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2825 )
         );
    snl_oa222x1 \ALUSHT/SHT/U569  ( .Z(\ALUSHT/SHT/n2575 ), .A(
        \ALUSHT/SHT/n2576 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2535 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2577 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_nand04x0 \ALUSHT/SHT/U659  ( .ZN(\ALUSHT/SHT/n2713 ), .A(
        \ALUSHT/SHT/n2603 ), .B(\ALUSHT/SHT/n2604 ), .C(\ALUSHT/SHT/n2605 ), 
        .D(\ALUSHT/SHT/n2606 ) );
    snl_oa2222x1 \ALUSHT/SHT/U765  ( .Z(\ALUSHT/SHT/n2580 ), .A(
        \ALUSHT/SHT/n2401 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2400 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2526 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2921 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi012x1 \ALUSHT/SHT/U827  ( .ZN(\ALUSHT/SHT/n2968 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[22] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_nand02x1 \ALUSHT/SHT/U469  ( .ZN(\ALUSHT/pkshtout[3] ), .A(
        \ALUSHT/SHT/n2309 ), .B(\ALUSHT/SHT/n2310 ) );
    snl_nand02x1 \ALUSHT/SHT/U472  ( .ZN(\ALUSHT/pkshtout[6] ), .A(
        \ALUSHT/SHT/n2315 ), .B(\ALUSHT/SHT/n2316 ) );
    snl_oai012x1 \ALUSHT/SHT/U800  ( .ZN(\ALUSHT/SHT/n2945 ), .A(
        \ALUSHT/SHT/n2522 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_invx05 \ALUSHT/SHT/U990  ( .ZN(\ALUSHT/SHT/n3071 ), .A(
        \ALUSHT/SHT/n2439 ) );
    snl_invx05 \ALUSHT/SHT/U742  ( .ZN(\ALUSHT/SHT/n2478 ), .A(
        \ALUSHT/SHT/n2379 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U759  ( .ZN(\ALUSHT/SHT/n2927 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[25] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[26] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[27] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[24] ) );
    snl_aoi022x1 \ALUSHT/SHT/U1097  ( .ZN(\ALUSHT/SHT/n2800 ), .A(
        \ALUSHT/SHT/n2611 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n3085 ), 
        .D(\phshtd[4] ) );
    snl_invx05 \ALUSHT/SHT/U1107  ( .ZN(\ALUSHT/SHT/n3092 ), .A(
        \ALUSHT/SHT/n2993 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U281  ( .ZN(\ALUSHT/SHT/n2526 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[11] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[12] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[13] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[10] ) );
    snl_aoi022x1 \ALUSHT/SHT/U311  ( .ZN(\ALUSHT/SHT/n2654 ), .A(
        \pgaluina[15] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[14] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi222x0 \ALUSHT/SHT/U336  ( .ZN(\ALUSHT/SHT/n2303 ), .A(
        \ALUSHT/SHT/n2645 ), .B(\pgaluina[0] ), .C(\ALUSHT/SHT/n2644 ), .D(
        \pgaluina[24] ), .E(\ALUSHT/SHT/n2635 ), .F(\ALUSHT/SHT/n2908 ) );
    snl_aoi122x0 \ALUSHT/SHT/U343  ( .ZN(\ALUSHT/SHT/n2339 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[10] ), .C(\pgaluina[18] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi122x0 \ALUSHT/SHT/U344  ( .ZN(\ALUSHT/SHT/n2337 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[9] ), .C(\pgaluina[17] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U363  ( .ZN(\ALUSHT/SHT/n2306 ), .A(
        \ALUSHT/SHT/n2450 ), .B(\ALUSHT/SHT/n2721 ), .C(\ALUSHT/SHT/n2461 ), 
        .D(\ALUSHT/SHT/n2723 ), .E(\pgaluina[9] ), .F(\ALUSHT/SHT/n2634 ), .G(
        \ALUSHT/SHT/n2690 ), .H(\ALUSHT/SHT/n2639 ) );
    snl_oai2222x0 \ALUSHT/SHT/U642  ( .ZN(\ALUSHT/SHT/n2479 ), .A(
        \ALUSHT/SHT/n2671 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2672 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2673 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2674 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_invx05 \ALUSHT/SHT/U1120  ( .ZN(\ALUSHT/SHT/n2992 ), .A(
        \ALUSHT/SHT/n2990 ) );
    snl_oai2222x0 \ALUSHT/SHT/U890  ( .ZN(\ALUSHT/SHT/n2877 ), .A(
        \ALUSHT/SHT/n2934 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2938 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2933 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2932 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai2222x0 \ALUSHT/SHT/U900  ( .ZN(\ALUSHT/SHT/n2735 ), .A(
        \ALUSHT/SHT/n3028 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2991 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2996 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3001 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oa022x1 \ALUSHT/SHT/U555  ( .Z(\ALUSHT/SHT/n2533 ), .A(
        \ALUSHT/SHT/n2523 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2393 ), 
        .D(\ALUSHT/SHT/n2399 ) );
    snl_aoi222x0 \ALUSHT/SHT/U572  ( .ZN(\ALUSHT/SHT/n2583 ), .A(
        \ALUSHT/SHT/n2584 ), .B(\ALUSHT/SHT/n2498 ), .C(\ALUSHT/SHT/n2530 ), 
        .D(\ALUSHT/SHT/n2537 ), .E(\ALUSHT/SHT/n2585 ), .F(\ALUSHT/SHT/n2503 )
         );
    snl_invx05 \ALUSHT/SHT/U927  ( .ZN(\ALUSHT/SHT/n3043 ), .A(
        \ALUSHT/SHT/n2887 ) );
    snl_invx1 \ALUSHT/SHT/U381  ( .ZN(\ALUSHT/SHT/n2390 ), .A(
        \ALUSHT/SHT/n2388 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U386  ( .ZN(\ALUSHT/SHT/n2325 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2895 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2901 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[19] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[11] ) );
    snl_aoi123x2 \ALUSHT/SHT/U407  ( .ZN(\ALUSHT/SHT/n2371 ), .A(
        \ALUSHT/SHT/n2379 ), .B(\ALUSHT/SHT/n2380 ), .C(exetype1), .D(
        \phshtd[5] ), .E(\ALUSHT/SHT/n2377 ), .F(\ALUSHT/SHT/n2378 ) );
    snl_aoi222x2 \ALUSHT/SHT/U420  ( .ZN(\ALUSHT/SHT/n2587 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[30] ), .C(\ALUSHT/SHT/n2505 ), .D(
        \pgaluina[29] ), .E(\ALUSHT/SHT/n2500 ), .F(\pgaluina[31] ) );
    snl_nand04x0 \ALUSHT/SHT/U665  ( .ZN(\ALUSHT/SHT/n2719 ), .A(
        \ALUSHT/SHT/n2553 ), .B(\ALUSHT/SHT/n2556 ), .C(\ALUSHT/SHT/n2560 ), 
        .D(\ALUSHT/SHT/n2563 ) );
    snl_aoi012x1 \ALUSHT/SHT/U852  ( .ZN(\ALUSHT/SHT/n2998 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[25] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_aoi122x0 \ALUSHT/SHT/U949  ( .ZN(\ALUSHT/SHT/n2689 ), .A(
        \ALUSHT/SHT/n2975 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n2973 ), 
        .D(\ALUSHT/SHT/n2298 ), .E(\ALUSHT/SHT/n2747 ) );
    snl_nand02x1 \ALUSHT/SHT/U1055  ( .ZN(\ALUSHT/SHT/n2858 ), .A(
        \ALUSHT/SHT/n2856 ), .B(\ALUSHT/SHT/n2855 ) );
    snl_oai122x0 \ALUSHT/SHT/U1072  ( .ZN(\ALUSHT/SHT/n2891 ), .A(
        \ALUSHT/SHT/n3041 ), .B(\ALUSHT/SHT/n2536 ), .C(\ALUSHT/SHT/n3085 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2886 ) );
    snl_nand02x1 \ALUSHT/SHT/U597  ( .ZN(\ALUSHT/SHT/n2621 ), .A(exetype1), 
        .B(\ALUSHT/SHT/n2622 ) );
    snl_aoi222x0 \ALUSHT/SHT/U680  ( .ZN(\ALUSHT/SHT/n2789 ), .A(
        \ALUSHT/SHT/n2437 ), .B(\ALUSHT/SHT/n2790 ), .C(\ALUSHT/SHT/n2791 ), 
        .D(\ALUSHT/SHT/n2792 ), .E(\ALUSHT/SHT/n2480 ), .F(\ALUSHT/SHT/n2793 )
         );
    snl_invx05 \ALUSHT/SHT/U710  ( .ZN(\ALUSHT/SHT/n2694 ), .A(
        \ALUSHT/SHT/n2402 ) );
    snl_invx05 \ALUSHT/SHT/U737  ( .ZN(\ALUSHT/SHT/n2915 ), .A(
        \ALUSHT/SHT/n2413 ) );
    snl_oai2222x0 \ALUSHT/SHT/U875  ( .ZN(\ALUSHT/SHT/n2829 ), .A(
        \ALUSHT/SHT/n3010 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n3013 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3012 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3011 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_aoi122x0 \ALUSHT/SHT/U969  ( .ZN(\ALUSHT/SHT/n3061 ), .A(
        \pgaluina[17] ), .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(
        \ALUSHT/SHT/n2999 ), .E(\ALUSHT/SHT/n2419 ) );
    snl_oai222x0 \ALUSHT/SHT/U1075  ( .ZN(\ALUSHT/SHT/n2888 ), .A(
        \ALUSHT/SHT/n3042 ), .B(\ALUSHT/SHT/n2638 ), .C(\phshtd[4] ), .D(
        \ALUSHT/SHT/n2474 ), .E(\ALUSHT/SHT/n3041 ), .F(\ALUSHT/SHT/n2640 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1052  ( .ZN(\ALUSHT/SHT/n2851 ), .A(
        \ALUSHT/SHT/n3102 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3095 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3097 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3099 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nand02x2 \ALUSHT/SHT/U400  ( .ZN(\ALUSHT/SHT/n2510 ), .A(\phshtd[5] ), 
        .B(\ALUSHT/SHT/n2382 ) );
    snl_aoi122x2 \ALUSHT/SHT/U427  ( .ZN(\ALUSHT/SHT/n2363 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[6] ), .C(\pgaluina[30] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_oai012x1 \ALUSHT/SHT/U590  ( .ZN(\ALUSHT/SHT/n2610 ), .A(
        \ALUSHT/SHT/n2611 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2397 ) );
    snl_aoi222x0 \ALUSHT/SHT/U687  ( .ZN(\ALUSHT/SHT/n2352 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2832 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2833 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2827 )
         );
    snl_nor02x1 \ALUSHT/SHT/U730  ( .ZN(\ALUSHT/SHT/n2460 ), .A(
        \ALUSHT/SHT/n2640 ), .B(\ALUSHT/SHT/n2626 ) );
    snl_aoi022x1 \ALUSHT/SHT/U872  ( .ZN(\ALUSHT/SHT/n3011 ), .A(
        \pgaluina[22] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[21] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_invx05 \ALUSHT/SHT/U717  ( .ZN(\ALUSHT/SHT/n2849 ), .A(
        \ALUSHT/SHT/n2642 ) );
    snl_aoi222x1 \ALUSHT/SHT/U449  ( .ZN(\ALUSHT/SHT/n2838 ), .A(
        \ALUSHT/SHT/n2548 ), .B(\ALUSHT/SHT/n2839 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2785 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2783 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U779  ( .ZN(\ALUSHT/SHT/n2549 ), .A(
        \ALUSHT/SHT/n2925 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2528 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2385 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2529 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi012x1 \ALUSHT/SHT/U855  ( .ZN(\ALUSHT/SHT/n3000 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[17] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_nor04x0 \ALUSHT/SHT/U662  ( .ZN(\ALUSHT/SHT/n2716 ), .A(
        \ALUSHT/SHT/n2712 ), .B(\ALUSHT/SHT/n2713 ), .C(\ALUSHT/SHT/n2714 ), 
        .D(\ALUSHT/SHT/n2715 ) );
    snl_nand04x0 \ALUSHT/SHT/U1090  ( .ZN(\ALUSHT/SHT/n2666 ), .A(
        \ALUSHT/SHT/n2718 ), .B(\ALUSHT/SHT/n2717 ), .C(\ALUSHT/SHT/n2720 ), 
        .D(\ALUSHT/SHT/n2716 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1100  ( .ZN(\ALUSHT/SHT/n3111 ), .A(
        \ALUSHT/SHT/n2688 ), .B(\ALUSHT/SHT/n2504 ), .C(\ALUSHT/SHT/n2690 ), 
        .D(\phshtd[0] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U358  ( .ZN(\ALUSHT/SHT/n2309 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2754 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2763 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[27] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[3] ) );
    snl_ao222x1 \ALUSHT/SHT/U364  ( .Z(\ALUSHT/SHT/n2297 ), .A(
        \ALUSHT/SHT/n2656 ), .B(\ALUSHT/SHT/n2804 ), .C(\ALUSHT/SHT/n2805 ), 
        .D(\ALUSHT/SHT/n2441 ), .E(\ALUSHT/SHT/n2655 ), .F(\ALUSHT/SHT/n2806 )
         );
    snl_oai222x0 \ALUSHT/SHT/U552  ( .ZN(\ALUSHT/SHT/n2475 ), .A(
        \ALUSHT/SHT/n2525 ), .B(\ALUSHT/SHT/n2399 ), .C(\ALUSHT/SHT/n2395 ), 
        .D(\ALUSHT/SHT/n2402 ), .E(\ALUSHT/SHT/n2526 ), .F(\ALUSHT/SHT/n2392 )
         );
    snl_oai122x0 \ALUSHT/SHT/U575  ( .ZN(\ALUSHT/SHT/n2591 ), .A(
        \ALUSHT/SHT/n2592 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2593 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_oai2222x0 \ALUSHT/SHT/U920  ( .ZN(\ALUSHT/SHT/n2740 ), .A(
        \ALUSHT/SHT/n3040 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2976 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2980 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3018 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_aoi023x0 \ALUSHT/SHT/U645  ( .ZN(\ALUSHT/SHT/n2680 ), .A(
        \ALUSHT/SHT/n2681 ), .B(\ALUSHT/SHT/n2427 ), .C(\ALUSHT/SHT/n2435 ), 
        .D(\ALUSHT/SHT/n2682 ), .E(\ALUSHT/SHT/n2683 ) );
    snl_oai2222x0 \ALUSHT/SHT/U897  ( .ZN(\ALUSHT/SHT/n2734 ), .A(
        \ALUSHT/SHT/n2958 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3017 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n3026 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n2955 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_oai012x1 \ALUSHT/SHT/U907  ( .ZN(\ALUSHT/SHT/n2405 ), .A(
        \ALUSHT/SHT/n3003 ), .B(\ALUSHT/SHT/n2500 ), .C(\ALUSHT/SHT/n2540 ) );
    snl_aoi012x1 \ALUSHT/SHT/U1000  ( .ZN(\ALUSHT/SHT/n3077 ), .A(
        \ALUSHT/SHT/n3033 ), .B(\ALUSHT/SHT/n2390 ), .C(\ALUSHT/SHT/n2473 ) );
    snl_aoi223x1 \ALUSHT/SHT/U452  ( .ZN(\ALUSHT/SHT/n2860 ), .A(
        \ALUSHT/SHT/n2539 ), .B(\ALUSHT/SHT/n2792 ), .C(\ALUSHT/SHT/n2659 ), 
        .D(\ALUSHT/SHT/n2662 ), .E(\ALUSHT/SHT/n2793 ), .F(\ALUSHT/SHT/n2810 ), 
        .G(\ALUSHT/SHT/n2861 ) );
    snl_nand02x1 \ALUSHT/SHT/U475  ( .ZN(\ALUSHT/pkshtout[9] ), .A(
        \ALUSHT/SHT/n2321 ), .B(\ALUSHT/SHT/n2322 ) );
    snl_invx05 \ALUSHT/SHT/U549  ( .ZN(\ALUSHT/SHT/n2521 ), .A(\pgaluina[1] )
         );
    snl_aoi222x0 \ALUSHT/SHT/U679  ( .ZN(\ALUSHT/SHT/n2364 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2786 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2787 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2677 )
         );
    snl_nand02x1 \ALUSHT/SHT/U1027  ( .ZN(\ALUSHT/SHT/n2815 ), .A(
        \ALUSHT/SHT/n2813 ), .B(\ALUSHT/SHT/n2809 ) );
    snl_invx05 \ALUSHT/SHT/U745  ( .ZN(\ALUSHT/SHT/n2695 ), .A(
        \ALUSHT/SHT/n2918 ) );
    snl_oai012x1 \ALUSHT/SHT/U807  ( .ZN(\ALUSHT/SHT/n2775 ), .A(
        \ALUSHT/SHT/n2414 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_oai222x0 \ALUSHT/SHT/U997  ( .ZN(\ALUSHT/SHT/n2443 ), .A(
        \ALUSHT/SHT/n3019 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n3020 ), 
        .D(\ALUSHT/SHT/n2638 ), .E(\phshtd[4] ), .F(\ALUSHT/SHT/n2544 ) );
    snl_nand02x1 \ALUSHT/SHT/U527  ( .ZN(\ALUSHT/SHT/n2501 ), .A(
        \ALUSHT/SHT/n2382 ), .B(\ALUSHT/SHT/n2427 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U762  ( .ZN(\ALUSHT/SHT/n2929 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[17] ), .C(\pgaluina[18] ), .D(
        \ALUSHT/SHT/n2541 ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[19] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[16] ) );
    snl_invx05 \ALUSHT/SHT/U820  ( .ZN(\ALUSHT/SHT/n2652 ), .A(
        \ALUSHT/SHT/n2491 ) );
    snl_oai2222x0 \ALUSHT/SHT/U869  ( .ZN(\ALUSHT/SHT/n2872 ), .A(
        \ALUSHT/SHT/n3005 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n3008 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3007 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3006 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_and02x1 \ALUSHT/SHT/U617  ( .Z(\ALUSHT/SHT/n2641 ), .A(
        \ALUSHT/SHT/n2635 ), .B(\phshtd[0] ) );
    snl_oa012x1 \ALUSHT/SHT/U955  ( .Z(\ALUSHT/SHT/n3054 ), .A(\phshtd[2] ), 
        .B(\ALUSHT/SHT/n2558 ), .C(\ALUSHT/SHT/n2653 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1049  ( .ZN(\ALUSHT/SHT/n2845 ), .A(
        \ALUSHT/SHT/n3100 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3091 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3096 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3098 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nand02x1 \ALUSHT/SHT/U630  ( .ZN(\ALUSHT/SHT/n2657 ), .A(
        \ALUSHT/SHT/n2537 ), .B(\ALUSHT/SHT/n2298 ) );
    snl_oai012x1 \ALUSHT/SHT/U787  ( .ZN(\ALUSHT/SHT/n2935 ), .A(
        \ALUSHT/SHT/n2934 ), .B(\ALUSHT/SHT/n2500 ), .C(\ALUSHT/SHT/n2551 ) );
    snl_nand02x1 \ALUSHT/SHT/U490  ( .ZN(\ALUSHT/pkshtout[24] ), .A(
        \ALUSHT/SHT/n2351 ), .B(\ALUSHT/SHT/n2352 ) );
    snl_aoi012x1 \ALUSHT/SHT/U293  ( .ZN(\ALUSHT/SHT/n2737 ), .A(
        \ALUSHT/SHT/n2651 ), .B(\pgaluina[6] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oa2222x1 \ALUSHT/SHT/U324  ( .Z(\ALUSHT/SHT/n2570 ), .A(
        \ALUSHT/SHT/n2919 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2920 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2523 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2524 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi112x0 \ALUSHT/SHT/U500  ( .ZN(\ALUSHT/SHT/n2369 ), .A(\phshtd[5] ), 
        .B(\ALUSHT/SHT/n2377 ), .C(exetype1), .D(\ALUSHT/SHT/n2378 ) );
    snl_aoi222x0 \ALUSHT/SHT/U947  ( .ZN(\ALUSHT/SHT/n2466 ), .A(
        \ALUSHT/SHT/n2685 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2945 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2386 ), .F(\ALUSHT/SHT/n2687 )
         );
    snl_ao122x1 \ALUSHT/SHT/U972  ( .Z(\ALUSHT/SHT/n3063 ), .A(\pgaluina[19] ), 
        .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(\ALUSHT/SHT/n2995 ), 
        .E(\ALUSHT/SHT/n2419 ) );
    snl_invx05 \ALUSHT/SHT/U535  ( .ZN(\ALUSHT/SHT/n2509 ), .A(\pgaluina[14] )
         );
    snl_nand02x1 \ALUSHT/SHT/U605  ( .ZN(\ALUSHT/SHT/n2629 ), .A(
        \ALUSHT/SHT/n2506 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_invx05 \ALUSHT/SHT/U795  ( .ZN(\ALUSHT/SHT/n2942 ), .A(
        \ALUSHT/SHT/n2823 ) );
    snl_and02x1 \ALUSHT/SHT/U622  ( .Z(\ALUSHT/SHT/n2497 ), .A(
        \ALUSHT/SHT/n2650 ), .B(\ALUSHT/SHT/n2542 ) );
    snl_oai122x0 \ALUSHT/SHT/U960  ( .ZN(\ALUSHT/SHT/n2763 ), .A(
        \ALUSHT/SHT/n3052 ), .B(\ALUSHT/SHT/n2642 ), .C(\ALUSHT/SHT/n3053 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n2756 ) );
    snl_aoi122x0 \ALUSHT/SHT/U303  ( .ZN(\ALUSHT/SHT/n3046 ), .A(\pgaluina[5] 
        ), .B(\ALUSHT/SHT/n2459 ), .C(\ALUSHT/SHT/n2957 ), .D(
        \ALUSHT/SHT/n2298 ), .E(\ALUSHT/SHT/n2460 ) );
    snl_aoi112x0 \ALUSHT/SHT/U512  ( .ZN(\ALUSHT/SHT/n2422 ), .A(
        \ALUSHT/SHT/n2423 ), .B(\pgaluina[29] ), .C(\ALUSHT/SHT/n2424 ), .D(
        \ALUSHT/SHT/n2419 ) );
    snl_invx2 \ALUSHT/SHT/U388  ( .ZN(\ALUSHT/SHT/n2382 ), .A(\phshtd[4] ) );
    snl_nand02x1 \ALUSHT/SHT/U482  ( .ZN(\ALUSHT/pkshtout[16] ), .A(
        \ALUSHT/SHT/n2335 ), .B(\ALUSHT/SHT/n2336 ) );
    snl_aoi012x1 \ALUSHT/SHT/U599  ( .ZN(\ALUSHT/SHT/n2624 ), .A(
        \ALUSHT/SHT/n2370 ), .B(\ALUSHT/SHT/n2372 ), .C(\ALUSHT/SHT/n2623 ) );
    snl_invx05 \ALUSHT/SHT/U739  ( .ZN(\ALUSHT/SHT/n2432 ), .A(
        \ALUSHT/SHT/n2628 ) );
    snl_aoi222x1 \ALUSHT/SHT/U409  ( .ZN(\ALUSHT/SHT/n2856 ), .A(
        \ALUSHT/SHT/n2498 ), .B(\ALUSHT/SHT/n2857 ), .C(\ALUSHT/SHT/n2849 ), 
        .D(\ALUSHT/SHT/n2759 ), .E(\ALUSHT/SHT/n2548 ), .F(\ALUSHT/SHT/n2757 )
         );
    snl_nand02x1 \ALUSHT/SHT/U467  ( .ZN(\ALUSHT/pkshtout[1] ), .A(
        \ALUSHT/SHT/n2305 ), .B(\ALUSHT/SHT/n2306 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U757  ( .ZN(\ALUSHT/SHT/n2924 ), .A(
        \pgaluina[18] ), .B(\ALUSHT/SHT/n2631 ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[19] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[20] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[17] ) );
    snl_ao012x1 \ALUSHT/SHT/U815  ( .Z(\ALUSHT/SHT/n2458 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[9] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1099  ( .ZN(\ALUSHT/SHT/n2484 ), .A(
        \ALUSHT/SHT/n2684 ), .B(\ALUSHT/SHT/n2504 ), .C(\ALUSHT/SHT/n2462 ), 
        .D(\phshtd[0] ) );
    snl_invx05 \ALUSHT/SHT/U1109  ( .ZN(\ALUSHT/SHT/n3025 ), .A(
        \ALUSHT/SHT/n2948 ) );
    snl_nand04x0 \ALUSHT/SHT/U985  ( .ZN(\ALUSHT/SHT/n3069 ), .A(
        \ALUSHT/SHT/n2849 ), .B(\ALUSHT/SHT/n2435 ), .C(\ALUSHT/SHT/n2910 ), 
        .D(\pgaluina[30] ) );
    snl_oa2222x1 \ALUSHT/SHT/U277  ( .Z(\ALUSHT/SHT/n2593 ), .A(
        \ALUSHT/SHT/n2664 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2918 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2920 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2919 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U280  ( .ZN(\ALUSHT/SHT/n2524 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[12] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[13] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[14] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[11] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U288  ( .ZN(\ALUSHT/SHT/n2532 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[5] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[6] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[7] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[4] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U351  ( .ZN(\ALUSHT/SHT/n2317 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2730 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2736 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[31] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[7] ) );
    snl_aoi122x2 \ALUSHT/SHT/U440  ( .ZN(\ALUSHT/SHT/n2576 ), .A(
        \ALUSHT/SHT/n2931 ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2700 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2914 ) );
    snl_aoi012x1 \ALUSHT/SHT/U832  ( .ZN(\ALUSHT/SHT/n2977 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[26] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_invx05 \ALUSHT/SHT/U540  ( .ZN(\ALUSHT/SHT/n2514 ), .A(\pgaluina[10] )
         );
    snl_aoi222x0 \ALUSHT/SHT/U670  ( .ZN(\ALUSHT/SHT/n2748 ), .A(
        \ALUSHT/SHT/n2662 ), .B(\ALUSHT/SHT/n2749 ), .C(\ALUSHT/SHT/n2480 ), 
        .D(\ALUSHT/SHT/n2750 ), .E(\ALUSHT/SHT/n2437 ), .F(\ALUSHT/SHT/n2751 )
         );
    snl_oa122x1 \ALUSHT/SHT/U770  ( .Z(\ALUSHT/SHT/n2557 ), .A(
        \ALUSHT/SHT/n2928 ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2926 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2697 ) );
    snl_oai2222x0 \ALUSHT/SHT/U929  ( .ZN(\ALUSHT/SHT/n2843 ), .A(
        \ALUSHT/SHT/n2940 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2654 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2943 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2941 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_invx05 \ALUSHT/SHT/U1012  ( .ZN(\ALUSHT/SHT/n3083 ), .A(
        \ALUSHT/SHT/n2819 ) );
    snl_oai122x0 \ALUSHT/SHT/U1035  ( .ZN(\ALUSHT/SHT/n2826 ), .A(
        \ALUSHT/SHT/n2580 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2937 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2822 ) );
    snl_aoi222x0 \ALUSHT/SHT/U932  ( .ZN(\ALUSHT/SHT/n3047 ), .A(
        \ALUSHT/SHT/n2458 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2956 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2386 ), .F(\ALUSHT/SHT/n3048 )
         );
    snl_invx1 \ALUSHT/SHT/U376  ( .ZN(\ALUSHT/SHT/n2686 ), .A(
        \ALUSHT/SHT/n2614 ) );
    snl_oai2222x0 \ALUSHT/SHT/U885  ( .ZN(\ALUSHT/SHT/n2765 ), .A(
        \ALUSHT/SHT/n2654 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2667 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2617 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2618 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1009  ( .ZN(\ALUSHT/SHT/n2790 ), .A(
        \ALUSHT/SHT/n3008 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n3012 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3011 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3010 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai2222x0 \ALUSHT/SHT/U915  ( .ZN(\ALUSHT/SHT/n2741 ), .A(
        \ALUSHT/SHT/n3034 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3031 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n3029 ), .F(\ALUSHT/SHT/n2642 ), 
        .G(\ALUSHT/SHT/n3035 ), .H(\ALUSHT/SHT/n2454 ) );
    snl_invx1 \ALUSHT/SHT/U393  ( .ZN(\ALUSHT/SHT/n2504 ), .A(\phshtd[0] ) );
    snl_oai222x0 \ALUSHT/SHT/U567  ( .ZN(\ALUSHT/SHT/n2567 ), .A(
        \ALUSHT/SHT/n2568 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2569 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2570 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_oai122x0 \ALUSHT/SHT/U582  ( .ZN(\ALUSHT/SHT/n2602 ), .A(
        \ALUSHT/SHT/n2566 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2564 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_nor04x0 \ALUSHT/SHT/U657  ( .ZN(\ALUSHT/SHT/n2711 ), .A(
        \ALUSHT/SHT/n2710 ), .B(\ALUSHT/SHT/n2604 ), .C(\ALUSHT/SHT/n2608 ), 
        .D(\ALUSHT/SHT/n2609 ) );
    snl_oai122x0 \ALUSHT/SHT/U829  ( .ZN(\ALUSHT/SHT/n2973 ), .A(
        \ALUSHT/SHT/n2512 ), .B(\ALUSHT/SHT/n2413 ), .C(\ALUSHT/SHT/n2972 ), 
        .D(\ALUSHT/SHT/n2382 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_invx05 \ALUSHT/SHT/U860  ( .ZN(\ALUSHT/SHT/n3002 ), .A(
        \ALUSHT/SHT/n2479 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1082  ( .ZN(\ALUSHT/SHT/n2899 ), .A(
        \ALUSHT/SHT/n3109 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n2947 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n2950 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3108 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_invx05 \ALUSHT/SHT/U1112  ( .ZN(\ALUSHT/SHT/n2936 ), .A(
        \ALUSHT/SHT/n2935 ) );
    snl_aoi222x2 \ALUSHT/SHT/U412  ( .ZN(\ALUSHT/SHT/n2862 ), .A(
        \ALUSHT/SHT/n2498 ), .B(\ALUSHT/SHT/n2863 ), .C(\ALUSHT/SHT/n2849 ), 
        .D(\ALUSHT/SHT/n2790 ), .E(\ALUSHT/SHT/n2548 ), .F(\ALUSHT/SHT/n2819 )
         );
    snl_aoi122x2 \ALUSHT/SHT/U435  ( .ZN(\ALUSHT/SHT/n2568 ), .A(
        \ALUSHT/SHT/n2389 ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2695 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2914 ) );
    snl_aoi222x0 \ALUSHT/SHT/U695  ( .ZN(\ALUSHT/SHT/n2338 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2869 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2870 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2865 )
         );
    snl_invx05 \ALUSHT/SHT/U705  ( .ZN(\ALUSHT/SHT/n2503 ), .A(
        \ALUSHT/SHT/n2502 ) );
    snl_invx05 \ALUSHT/SHT/U722  ( .ZN(\ALUSHT/SHT/n2437 ), .A(
        \ALUSHT/SHT/n2451 ) );
    snl_aoi012x1 \ALUSHT/SHT/U847  ( .ZN(\ALUSHT/SHT/n2993 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[27] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1067  ( .ZN(\ALUSHT/SHT/n2878 ), .A(
        \ALUSHT/SHT/n2986 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3100 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3103 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3106 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_invx1 \ALUSHT/SHT/U318  ( .ZN(\ALUSHT/SHT/n2910 ), .A(
        \ALUSHT/SHT/n2612 ) );
    snl_oai122x0 \ALUSHT/SHT/U509  ( .ZN(\ALUSHT/SHT/n2411 ), .A(
        \ALUSHT/SHT/n2382 ), .B(\ALUSHT/SHT/n2412 ), .C(\ALUSHT/SHT/n2413 ), 
        .D(\ALUSHT/SHT/n2414 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_aoi222x0 \ALUSHT/SHT/U337  ( .ZN(\ALUSHT/SHT/n2368 ), .A(
        \ALUSHT/SHT/n2635 ), .B(\ALUSHT/SHT/n2780 ), .C(\ALUSHT/SHT/n2781 ), 
        .D(\ALUSHT/SHT/n2381 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[7] ) );
    snl_nor03x0 \ALUSHT/SHT/U499  ( .ZN(\ALUSHT/slaovf ), .A(
        \ALUSHT/SHT/n2375 ), .B(pkshterr), .C(\ALUSHT/SHT/n2376 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U639  ( .ZN(\ALUSHT/SHT/n2664 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[28] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[29] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[30] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[27] ) );
    snl_aoi022x1 \ALUSHT/SHT/U868  ( .ZN(\ALUSHT/SHT/n3008 ), .A(
        \pgaluina[26] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[25] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1040  ( .ZN(\ALUSHT/SHT/n2833 ), .A(
        \ALUSHT/SHT/n3097 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3078 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3088 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3095 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oa2222x1 \ALUSHT/SHT/U1048  ( .Z(\ALUSHT/SHT/n3100 ), .A(
        \ALUSHT/SHT/n3101 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2987 ), 
        .D(\ALUSHT/SHT/n2627 ), .E(\ALUSHT/SHT/n2990 ), .F(\ALUSHT/SHT/n2501 ), 
        .G(\ALUSHT/SHT/n2770 ), .H(\ALUSHT/SHT/n2638 ) );
    snl_oa012x1 \ALUSHT/SHT/U501  ( .Z(\ALUSHT/SHT/n2373 ), .A(
        \ALUSHT/SHT/n2381 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n2377 ) );
    snl_nand02x1 \ALUSHT/SHT/U526  ( .ZN(\ALUSHT/SHT/n2455 ), .A(
        \ALUSHT/SHT/n2498 ), .B(\ALUSHT/SHT/n2427 ) );
    snl_and02x1 \ALUSHT/SHT/U616  ( .Z(\ALUSHT/SHT/n2639 ), .A(
        \ALUSHT/SHT/n2635 ), .B(\ALUSHT/SHT/n2504 ) );
    snl_aoi022x1 \ALUSHT/SHT/U786  ( .ZN(\ALUSHT/SHT/n2934 ), .A(
        \pgaluina[31] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[30] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_invx05 \ALUSHT/SHT/U954  ( .ZN(\ALUSHT/SHT/n3053 ), .A(
        \ALUSHT/SHT/n2811 ) );
    snl_nor02x1 \ALUSHT/SHT/U631  ( .ZN(\ALUSHT/SHT/n2418 ), .A(
        \ALUSHT/SHT/n2374 ), .B(\ALUSHT/SHT/n2502 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U289  ( .ZN(\ALUSHT/SHT/n2393 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[4] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[5] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[6] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[3] ) );
    snl_aoi022x1 \ALUSHT/SHT/U310  ( .ZN(\ALUSHT/SHT/n2618 ), .A(
        \pgaluina[13] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[12] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_nand02x1 \ALUSHT/SHT/U491  ( .ZN(\ALUSHT/pkshtout[25] ), .A(
        \ALUSHT/SHT/n2353 ), .B(\ALUSHT/SHT/n2354 ) );
    snl_aoi023x0 \ALUSHT/SHT/U319  ( .ZN(\ALUSHT/SHT/n2442 ), .A(
        \ALUSHT/SHT/n2443 ), .B(\ALUSHT/SHT/n2441 ), .C(\ALUSHT/SHT/n2444 ), 
        .D(\ALUSHT/SHT/n2445 ), .E(\pgaluina[15] ) );
    snl_aoi122x0 \ALUSHT/SHT/U342  ( .ZN(\ALUSHT/SHT/n2341 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[11] ), .C(\pgaluina[19] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U359  ( .ZN(\ALUSHT/SHT/n2310 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2760 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2761 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[11] ), 
        .G(\ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2762 ) );
    snl_invx05 \ALUSHT/SHT/U548  ( .ZN(\ALUSHT/SHT/n2449 ), .A(\pgaluina[2] )
         );
    snl_aoi122x0 \ALUSHT/SHT/U973  ( .ZN(\ALUSHT/SHT/n3064 ), .A(
        \pgaluina[15] ), .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(
        \ALUSHT/SHT/n2982 ), .E(\ALUSHT/SHT/n2419 ) );
    snl_oai122x0 \ALUSHT/SHT/U1001  ( .ZN(\ALUSHT/SHT/n2786 ), .A(
        \ALUSHT/SHT/n3035 ), .B(\ALUSHT/SHT/n2657 ), .C(\ALUSHT/SHT/n3032 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n2782 ) );
    snl_invx05 \ALUSHT/SHT/U1026  ( .ZN(\ALUSHT/SHT/n2814 ), .A(
        \ALUSHT/SHT/n3090 ) );
    snl_aoi222x1 \ALUSHT/SHT/U448  ( .ZN(\ALUSHT/SHT/n2871 ), .A(
        \ALUSHT/SHT/n2662 ), .B(\ALUSHT/SHT/n2872 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2497 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2479 )
         );
    snl_aoi222x1 \ALUSHT/SHT/U453  ( .ZN(\ALUSHT/SHT/n2834 ), .A(
        \ALUSHT/SHT/n2548 ), .B(\ALUSHT/SHT/n2835 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2767 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2765 )
         );
    snl_nand02x1 \ALUSHT/SHT/U474  ( .ZN(\ALUSHT/pkshtout[8] ), .A(
        \ALUSHT/SHT/n2319 ), .B(\ALUSHT/SHT/n2320 ) );
    snl_aoi222x0 \ALUSHT/SHT/U678  ( .ZN(\ALUSHT/SHT/n2782 ), .A(
        \ALUSHT/SHT/n2656 ), .B(\ALUSHT/SHT/n2783 ), .C(\ALUSHT/SHT/n2784 ), 
        .D(\ALUSHT/SHT/n2441 ), .E(\ALUSHT/SHT/n2655 ), .F(\ALUSHT/SHT/n2785 )
         );
    snl_aoi2222x0 \ALUSHT/SHT/U744  ( .ZN(\ALUSHT/SHT/n2918 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[24] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[25] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[26] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[23] ) );
    snl_oai122x0 \ALUSHT/SHT/U806  ( .ZN(\ALUSHT/SHT/n2776 ), .A(
        \ALUSHT/SHT/n2517 ), .B(\ALUSHT/SHT/n2628 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n2948 ), .E(\ALUSHT/SHT/n2913 ) );
    snl_oai012x1 \ALUSHT/SHT/U996  ( .ZN(\ALUSHT/SHT/n2436 ), .A(
        \ALUSHT/SHT/n2509 ), .B(\ALUSHT/SHT/n2612 ), .C(\ALUSHT/SHT/n2626 ) );
    snl_oai2222x0 \ALUSHT/SHT/U763  ( .ZN(\ALUSHT/SHT/n2585 ), .A(
        \ALUSHT/SHT/n2927 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2928 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2930 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2929 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi012x1 \ALUSHT/SHT/U821  ( .ZN(\ALUSHT/SHT/n2961 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[24] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oai2222x0 \ALUSHT/SHT/U778  ( .ZN(\ALUSHT/SHT/n2547 ), .A(
        \ALUSHT/SHT/n2587 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2922 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2924 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2923 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_oa022x1 \ALUSHT/SHT/U553  ( .Z(\ALUSHT/SHT/n2527 ), .A(
        \ALUSHT/SHT/n2528 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2529 ), 
        .D(\ALUSHT/SHT/n2399 ) );
    snl_nor04x0 \ALUSHT/SHT/U663  ( .ZN(\ALUSHT/SHT/n2717 ), .A(
        \ALUSHT/SHT/n2589 ), .B(\ALUSHT/SHT/n2586 ), .C(\ALUSHT/SHT/n2583 ), 
        .D(\ALUSHT/SHT/n2581 ) );
    snl_invx05 \ALUSHT/SHT/U1091  ( .ZN(\ALUSHT/SHT/n2824 ), .A(
        \ALUSHT/SHT/n2493 ) );
    snl_invx05 \ALUSHT/SHT/U1101  ( .ZN(\ALUSHT/SHT/n2931 ), .A(
        \ALUSHT/SHT/n2587 ) );
    snl_aoi222x0 \ALUSHT/SHT/U365  ( .ZN(\ALUSHT/SHT/n3018 ), .A(
        \ALUSHT/SHT/n2488 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2960 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2489 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U921  ( .ZN(\ALUSHT/SHT/n2799 ), .A(
        \ALUSHT/SHT/n2618 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2670 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2667 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2617 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nand02x2 \ALUSHT/SHT/U380  ( .ZN(\ALUSHT/SHT/n2499 ), .A(
        \ALUSHT/SHT/n2386 ), .B(\ALUSHT/SHT/n2500 ) );
    snl_nand02x2 \ALUSHT/SHT/U401  ( .ZN(\ALUSHT/SHT/n2402 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n2386 ) );
    snl_aoi222x0 \ALUSHT/SHT/U574  ( .ZN(\ALUSHT/SHT/n2589 ), .A(
        \pgaluina[30] ), .B(\ALUSHT/SHT/n2498 ), .C(\ALUSHT/SHT/n2475 ), .D(
        \ALUSHT/SHT/n2537 ), .E(\ALUSHT/SHT/n2590 ), .F(\ALUSHT/SHT/n2503 ) );
    snl_nor02x1 \ALUSHT/SHT/U591  ( .ZN(\ALUSHT/SHT/n2445 ), .A(
        \ALUSHT/SHT/n2370 ), .B(\poshtfnc[0] ) );
    snl_oai222x0 \ALUSHT/SHT/U644  ( .ZN(\ALUSHT/SHT/n2677 ), .A(
        \ALUSHT/SHT/n2678 ), .B(\ALUSHT/SHT/n2619 ), .C(\ALUSHT/SHT/n2422 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\phshtd[1] ), .F(\ALUSHT/SHT/n2679 ) );
    snl_ao122x1 \ALUSHT/SHT/U896  ( .Z(\ALUSHT/SHT/n3024 ), .A(\pgaluina[7] ), 
        .B(\ALUSHT/SHT/n2459 ), .C(\ALUSHT/SHT/n3025 ), .D(\ALUSHT/SHT/n2298 ), 
        .E(\ALUSHT/SHT/n2460 ) );
    snl_invx05 \ALUSHT/SHT/U906  ( .ZN(\ALUSHT/SHT/n3031 ), .A(
        \ALUSHT/SHT/n2785 ) );
    snl_aoi222x0 \ALUSHT/SHT/U968  ( .ZN(\ALUSHT/SHT/n3060 ), .A(
        \ALUSHT/SHT/n3056 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2416 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2386 ), .F(\ALUSHT/SHT/n3058 )
         );
    snl_oai122x0 \ALUSHT/SHT/U1053  ( .ZN(\ALUSHT/SHT/n2854 ), .A(
        \ALUSHT/SHT/n2944 ), .B(\ALUSHT/SHT/n2454 ), .C(\ALUSHT/SHT/n2452 ), 
        .D(\ALUSHT/SHT/n2642 ), .E(\ALUSHT/SHT/n2852 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1074  ( .ZN(\ALUSHT/SHT/n2890 ), .A(
        \ALUSHT/SHT/n2991 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3103 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3106 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2986 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nor02x2 \ALUSHT/SHT/U392  ( .ZN(\ALUSHT/SHT/n2505 ), .A(
        \ALUSHT/SHT/n2500 ), .B(\ALUSHT/SHT/n2504 ) );
    snl_aoi222x1 \ALUSHT/SHT/U413  ( .ZN(\ALUSHT/SHT/n2813 ), .A(
        \ALUSHT/SHT/n2503 ), .B(\ALUSHT/SHT/n2814 ), .C(\ALUSHT/SHT/n2548 ), 
        .D(\ALUSHT/SHT/n2759 ), .E(\ALUSHT/SHT/n2498 ), .F(\ALUSHT/SHT/n2585 )
         );
    snl_aoi122x2 \ALUSHT/SHT/U426  ( .ZN(\ALUSHT/SHT/n2353 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[1] ), .C(\pgaluina[25] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi222x0 \ALUSHT/SHT/U686  ( .ZN(\ALUSHT/SHT/n2354 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2826 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2827 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2821 )
         );
    snl_invx05 \ALUSHT/SHT/U716  ( .ZN(\ALUSHT/SHT/n2548 ), .A(
        \ALUSHT/SHT/n2536 ) );
    snl_nor02x1 \ALUSHT/SHT/U731  ( .ZN(\ALUSHT/SHT/n2914 ), .A(
        \ALUSHT/SHT/n2366 ), .B(\ALUSHT/SHT/n2298 ) );
    snl_aoi022x1 \ALUSHT/SHT/U873  ( .ZN(\ALUSHT/SHT/n3012 ), .A(
        \pgaluina[20] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[19] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_oai012x1 \ALUSHT/SHT/U854  ( .ZN(\ALUSHT/SHT/n2999 ), .A(
        \ALUSHT/SHT/n2521 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U861  ( .ZN(\ALUSHT/SHT/n3003 ), .A(
        \pgaluina[15] ), .B(\ALUSHT/SHT/n2910 ), .C(\ALUSHT/SHT/n2917 ) );
    snl_aoi222x2 \ALUSHT/SHT/U434  ( .ZN(\ALUSHT/SHT/n3109 ), .A(
        \ALUSHT/SHT/n2957 ), .B(\ALUSHT/SHT/n2539 ), .C(\ALUSHT/SHT/n2431 ), 
        .D(\ALUSHT/SHT/n2694 ), .E(\ALUSHT/SHT/n3072 ), .F(\phshtd[2] ) );
    snl_oai122x0 \ALUSHT/SHT/U583  ( .ZN(\ALUSHT/SHT/n2603 ), .A(
        \ALUSHT/SHT/n2570 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2568 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi222x0 \ALUSHT/SHT/U694  ( .ZN(\ALUSHT/SHT/n2340 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2864 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2865 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2859 )
         );
    snl_invx05 \ALUSHT/SHT/U723  ( .ZN(\ALUSHT/SHT/n2723 ), .A(
        \ALUSHT/SHT/n2632 ) );
    snl_nor02x1 \ALUSHT/SHT/U704  ( .ZN(\ALUSHT/SHT/n2419 ), .A(
        \ALUSHT/SHT/n2637 ), .B(\ALUSHT/SHT/n2502 ) );
    snl_aoi222x0 \ALUSHT/SHT/U846  ( .ZN(\ALUSHT/SHT/n2991 ), .A(
        \ALUSHT/SHT/n2992 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2989 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2988 )
         );
    snl_oai222x0 \ALUSHT/SHT/U498  ( .ZN(pkshterr), .A(\ALUSHT/SHT/n2369 ), 
        .B(\ALUSHT/SHT/n2370 ), .C(\ALUSHT/SHT/n2371 ), .D(\ALUSHT/SHT/n2372 ), 
        .E(\ALUSHT/SHT/n2373 ), .F(\ALUSHT/SHT/n2374 ) );
    snl_ao012x1 \ALUSHT/SHT/U508  ( .Z(\ALUSHT/SHT/n2408 ), .A(\pgaluina[3] ), 
        .B(\ALUSHT/SHT/n2409 ), .C(\ALUSHT/SHT/n2410 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U350  ( .ZN(\ALUSHT/SHT/n2320 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2728 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2729 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[0] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2730 ) );
    snl_nand03x0 \ALUSHT/SHT/U638  ( .ZN(\ALUSHT/SHT/n2377 ), .A(
        \ALUSHT/SHT/n2661 ), .B(\ALUSHT/SHT/n2504 ), .C(\ALUSHT/SHT/n2663 ) );
    snl_oai122x0 \ALUSHT/SHT/U1066  ( .ZN(\ALUSHT/SHT/n2879 ), .A(
        \ALUSHT/SHT/n3019 ), .B(\ALUSHT/SHT/n2536 ), .C(\ALUSHT/SHT/n2544 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2876 ) );
    snl_aoi222x0 \ALUSHT/SHT/U671  ( .ZN(\ALUSHT/SHT/n2756 ), .A(
        \ALUSHT/SHT/n2662 ), .B(\ALUSHT/SHT/n2757 ), .C(\ALUSHT/SHT/n2480 ), 
        .D(\ALUSHT/SHT/n2758 ), .E(\ALUSHT/SHT/n2437 ), .F(\ALUSHT/SHT/n2759 )
         );
    snl_oai122x0 \ALUSHT/SHT/U1041  ( .ZN(\ALUSHT/SHT/n2836 ), .A(
        \ALUSHT/SHT/n2574 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3022 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2834 ) );
    snl_oai2222x0 \ALUSHT/SHT/U933  ( .ZN(\ALUSHT/SHT/n2744 ), .A(
        \ALUSHT/SHT/n3026 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3038 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n3047 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3017 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_nand02x2 \ALUSHT/SHT/U377  ( .ZN(\ALUSHT/SHT/n2614 ), .A(\phshtd[2] ), 
        .B(\ALUSHT/SHT/n2500 ) );
    snl_invx05 \ALUSHT/SHT/U541  ( .ZN(\ALUSHT/SHT/n2515 ), .A(\pgaluina[9] )
         );
    snl_oai222x0 \ALUSHT/SHT/U566  ( .ZN(\ALUSHT/SHT/n2563 ), .A(
        \ALUSHT/SHT/n2564 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2565 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2566 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U884  ( .ZN(\ALUSHT/SHT/n2730 ), .A(
        \ALUSHT/SHT/n3018 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2969 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2976 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2980 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_invx05 \ALUSHT/SHT/U914  ( .ZN(\ALUSHT/SHT/n3035 ), .A(
        \ALUSHT/SHT/n2839 ) );
    snl_or04x1 \ALUSHT/SHT/U656  ( .Z(\ALUSHT/SHT/n2710 ), .A(
        \ALUSHT/SHT/n2607 ), .B(\ALUSHT/SHT/n2606 ), .C(\ALUSHT/SHT/n2605 ), 
        .D(\ALUSHT/SHT/n2610 ) );
    snl_oai222x0 \ALUSHT/SHT/U1008  ( .ZN(\ALUSHT/SHT/n2793 ), .A(
        \ALUSHT/SHT/n3007 ), .B(\ALUSHT/SHT/n2615 ), .C(\ALUSHT/SHT/n3006 ), 
        .D(\ALUSHT/SHT/n2614 ), .E(\phshtd[2] ), .F(\ALUSHT/SHT/n3081 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U756  ( .ZN(\ALUSHT/SHT/n2923 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[22] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[23] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[24] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[21] ) );
    snl_aoi012x1 \ALUSHT/SHT/U828  ( .ZN(\ALUSHT/SHT/n2972 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[28] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1083  ( .ZN(\ALUSHT/SHT/n2900 ), .A(
        \ALUSHT/SHT/n2996 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3106 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2986 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2991 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_invx05 \ALUSHT/SHT/U1113  ( .ZN(\ALUSHT/SHT/n3101 ), .A(
        \ALUSHT/SHT/n2989 ) );
    snl_ao012x1 \ALUSHT/SHT/U814  ( .Z(\ALUSHT/SHT/n2957 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[13] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_oai012x1 \ALUSHT/SHT/U984  ( .ZN(\ALUSHT/SHT/n2429 ), .A(
        \ALUSHT/SHT/n2509 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U279  ( .ZN(\ALUSHT/SHT/n2930 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[13] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[14] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[15] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[12] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U292  ( .ZN(\ALUSHT/SHT/n2558 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[1] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[2] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[3] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[0] ) );
    snl_aoi122x0 \ALUSHT/SHT/U302  ( .ZN(\ALUSHT/SHT/n2457 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n2458 ), .C(\ALUSHT/SHT/n2459 ), 
        .D(\pgaluina[1] ), .E(\ALUSHT/SHT/n2460 ) );
    snl_oa2222x1 \ALUSHT/SHT/U325  ( .Z(\ALUSHT/SHT/n2566 ), .A(
        \ALUSHT/SHT/n2400 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2921 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2525 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2526 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi222x2 \ALUSHT/SHT/U441  ( .ZN(\ALUSHT/SHT/n2950 ), .A(
        \ALUSHT/SHT/n2949 ), .B(\ALUSHT/SHT/n2539 ), .C(\ALUSHT/SHT/n2775 ), 
        .D(\ALUSHT/SHT/n2694 ), .E(\ALUSHT/SHT/n2776 ), .F(\phshtd[2] ) );
    snl_nand02x1 \ALUSHT/SHT/U466  ( .ZN(\ALUSHT/pkshtout[0] ), .A(
        \ALUSHT/SHT/n2303 ), .B(\ALUSHT/SHT/n2304 ) );
    snl_oai122x0 \ALUSHT/SHT/U833  ( .ZN(\ALUSHT/SHT/n2978 ), .A(
        \ALUSHT/SHT/n2514 ), .B(\ALUSHT/SHT/n2413 ), .C(\ALUSHT/SHT/n2977 ), 
        .D(\ALUSHT/SHT/n2382 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1098  ( .ZN(\ALUSHT/SHT/n2805 ), .A(
        \ALUSHT/SHT/n2588 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n3087 ), 
        .D(\phshtd[4] ) );
    snl_invx05 \ALUSHT/SHT/U1108  ( .ZN(\ALUSHT/SHT/n2964 ), .A(
        \ALUSHT/SHT/n2960 ) );
    snl_nand02x1 \ALUSHT/SHT/U534  ( .ZN(\ALUSHT/SHT/n2508 ), .A(\phshtd[1] ), 
        .B(\ALUSHT/SHT/n2504 ) );
    snl_oai2222x0 \ALUSHT/SHT/U771  ( .ZN(\ALUSHT/SHT/n2857 ), .A(
        \ALUSHT/SHT/n2929 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2930 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2532 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2531 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi122x0 \ALUSHT/SHT/U928  ( .ZN(\ALUSHT/SHT/n3044 ), .A(
        \ALUSHT/SHT/n2935 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2887 ), 
        .D(\ALUSHT/SHT/n2298 ), .E(\ALUSHT/SHT/n2394 ) );
    snl_oai122x0 \ALUSHT/SHT/U1013  ( .ZN(\ALUSHT/SHT/n2797 ), .A(
        \ALUSHT/SHT/n3083 ), .B(\ALUSHT/SHT/n2454 ), .C(\ALUSHT/SHT/n3079 ), 
        .D(\ALUSHT/SHT/n2642 ), .E(\ALUSHT/SHT/n2789 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1034  ( .ZN(\ALUSHT/SHT/n2821 ), .A(
        \ALUSHT/SHT/n3095 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n3059 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3078 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3088 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_ao122x1 \ALUSHT/SHT/U946  ( .Z(\ALUSHT/SHT/n2687 ), .A(\pgaluina[4] ), 
        .B(\ALUSHT/SHT/n2459 ), .C(\ALUSHT/SHT/n2946 ), .D(\ALUSHT/SHT/n2298 ), 
        .E(\ALUSHT/SHT/n2460 ) );
    snl_nand02x1 \ALUSHT/SHT/U483  ( .ZN(\ALUSHT/pkshtout[17] ), .A(
        \ALUSHT/SHT/n2337 ), .B(\ALUSHT/SHT/n2338 ) );
    snl_nand02x1 \ALUSHT/SHT/U604  ( .ZN(\ALUSHT/SHT/n2465 ), .A(
        \ALUSHT/SHT/n2505 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_and02x1 \ALUSHT/SHT/U623  ( .Z(\ALUSHT/SHT/n2459 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\ALUSHT/SHT/n2427 ) );
    snl_oai2222x0 \ALUSHT/SHT/U794  ( .ZN(\ALUSHT/SHT/n2823 ), .A(
        \ALUSHT/SHT/n2938 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2941 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2940 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2939 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai2222x0 \ALUSHT/SHT/U961  ( .ZN(\ALUSHT/SHT/n2761 ), .A(
        \ALUSHT/SHT/n3047 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n2466 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n3055 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3038 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_aoi122x0 \ALUSHT/SHT/U513  ( .ZN(\ALUSHT/SHT/n2425 ), .A(
        \ALUSHT/SHT/n2426 ), .B(\ALUSHT/SHT/n2427 ), .C(\ALUSHT/SHT/n2428 ), 
        .D(\ALUSHT/SHT/n2429 ), .E(\ALUSHT/SHT/n2419 ) );
    snl_nor02x2 \ALUSHT/SHT/U295  ( .ZN(\ALUSHT/SHT/n2506 ), .A(\phshtd[0] ), 
        .B(\phshtd[1] ) );
    snl_invx1 \ALUSHT/SHT/U389  ( .ZN(\ALUSHT/SHT/n2428 ), .A(
        \ALUSHT/SHT/n2627 ) );
    snl_aoi222x2 \ALUSHT/SHT/U408  ( .ZN(\ALUSHT/SHT/n2905 ), .A(
        \ALUSHT/SHT/n2437 ), .B(\ALUSHT/SHT/n2829 ), .C(\ALUSHT/SHT/n2497 ), 
        .D(\ALUSHT/SHT/n2548 ), .E(\ALUSHT/SHT/n2480 ), .F(\ALUSHT/SHT/n2872 )
         );
    snl_nand02x1 \ALUSHT/SHT/U738  ( .ZN(\ALUSHT/SHT/n2916 ), .A(
        \ALUSHT/SHT/n2483 ), .B(\ALUSHT/SHT/n2382 ) );
    snl_invx05 \ALUSHT/SHT/U598  ( .ZN(\ALUSHT/SHT/n2623 ), .A(\poshtfnc[0] )
         );
    snl_aoi022x1 \ALUSHT/SHT/U305  ( .ZN(\ALUSHT/SHT/n2670 ), .A(\pgaluina[7] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[6] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_ao122x1 \ALUSHT/SHT/U514  ( .Z(\ALUSHT/SHT/n2430 ), .A(
        \ALUSHT/SHT/n2431 ), .B(\ALUSHT/SHT/n2427 ), .C(\ALUSHT/SHT/n2432 ), 
        .D(\pgaluina[13] ), .E(\ALUSHT/SHT/n2433 ) );
    snl_oa2222x1 \ALUSHT/SHT/U322  ( .Z(\ALUSHT/SHT/n2577 ), .A(
        \ALUSHT/SHT/n2923 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2924 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2528 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2925 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_nand02x1 \ALUSHT/SHT/U484  ( .ZN(\ALUSHT/pkshtout[18] ), .A(
        \ALUSHT/SHT/n2339 ), .B(\ALUSHT/SHT/n2340 ) );
    snl_nand02x1 \ALUSHT/SHT/U603  ( .ZN(\ALUSHT/SHT/n2628 ), .A(
        \ALUSHT/SHT/n2428 ), .B(\ALUSHT/SHT/n2477 ) );
    snl_nor02x1 \ALUSHT/SHT/U624  ( .ZN(\ALUSHT/SHT/n2651 ), .A(
        \ALUSHT/SHT/n2501 ), .B(\ALUSHT/SHT/n2652 ) );
    snl_invx05 \ALUSHT/SHT/U966  ( .ZN(\ALUSHT/SHT/n3059 ), .A(
        \ALUSHT/SHT/n3058 ) );
    snl_aoi022x1 \ALUSHT/SHT/U793  ( .ZN(\ALUSHT/SHT/n2941 ), .A(
        \pgaluina[19] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[18] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi122x0 \ALUSHT/SHT/U339  ( .ZN(\ALUSHT/SHT/n2347 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[14] ), .C(\pgaluina[22] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U357  ( .ZN(\ALUSHT/SHT/n2311 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2745 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2755 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[28] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[4] ) );
    snl_invx1 \ALUSHT/SHT/U370  ( .ZN(\ALUSHT/SHT/n2299 ), .A(
        \ALUSHT/SHT/n2682 ) );
    snl_aoi122x2 \ALUSHT/SHT/U428  ( .ZN(\ALUSHT/SHT/n2357 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[3] ), .C(\pgaluina[27] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_nand02x1 \ALUSHT/SHT/U533  ( .ZN(\ALUSHT/SHT/n2507 ), .A(\phshtd[0] ), 
        .B(\ALUSHT/SHT/n2500 ) );
    snl_aoi222x0 \ALUSHT/SHT/U688  ( .ZN(\ALUSHT/SHT/n2350 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2836 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2837 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2833 )
         );
    snl_invx05 \ALUSHT/SHT/U718  ( .ZN(\ALUSHT/SHT/n2662 ), .A(
        \ALUSHT/SHT/n2454 ) );
    snl_oai222x0 \ALUSHT/SHT/U941  ( .ZN(\ALUSHT/SHT/n2752 ), .A(
        \ALUSHT/SHT/n3049 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n3051 ), 
        .D(\ALUSHT/SHT/n2455 ), .E(\ALUSHT/SHT/n3050 ), .F(\ALUSHT/SHT/n2454 )
         );
    snl_invx1 \ALUSHT/SHT/U446  ( .ZN(\ALUSHT/SHT/n2441 ), .A(\phshtd[5] ) );
    snl_oai2222x0 \ALUSHT/SHT/U776  ( .ZN(\ALUSHT/SHT/n2868 ), .A(
        \ALUSHT/SHT/n2921 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2526 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2395 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2525 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_nand02x2 \ALUSHT/SHT/U461  ( .ZN(\ALUSHT/SHT/n2640 ), .A(\phshtd[4] ), 
        .B(\ALUSHT/SHT/n2427 ) );
    snl_oai012x1 \ALUSHT/SHT/U834  ( .ZN(\ALUSHT/SHT/n2979 ), .A(
        \ALUSHT/SHT/n2449 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_nand04x0 \ALUSHT/SHT/U651  ( .ZN(\ALUSHT/SHT/n2705 ), .A(
        \ALUSHT/SHT/n2581 ), .B(\ALUSHT/SHT/n2578 ), .C(\ALUSHT/SHT/n2575 ), 
        .D(\ALUSHT/SHT/n2571 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U751  ( .ZN(\ALUSHT/SHT/n2401 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[23] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[24] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[25] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[22] ) );
    snl_oai012x1 \ALUSHT/SHT/U813  ( .ZN(\ALUSHT/SHT/n2956 ), .A(
        \ALUSHT/SHT/n2521 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_ao122x1 \ALUSHT/SHT/U983  ( .Z(\ALUSHT/SHT/n2426 ), .A(\pgaluina[22] ), 
        .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(\ALUSHT/SHT/n2967 ), 
        .E(\ALUSHT/SHT/n2419 ) );
    snl_oai122x0 \ALUSHT/SHT/U898  ( .ZN(\ALUSHT/SHT/n3027 ), .A(
        \ALUSHT/SHT/n2985 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2983 ), 
        .D(\ALUSHT/SHT/n2427 ), .E(\ALUSHT/SHT/n2732 ) );
    snl_oa222x1 \ALUSHT/SHT/U1033  ( .Z(\ALUSHT/SHT/n3095 ), .A(
        \ALUSHT/SHT/n3068 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2977 ), 
        .D(\ALUSHT/SHT/n2501 ), .E(\ALUSHT/SHT/n3067 ), .F(\ALUSHT/SHT/n2427 )
         );
    snl_oai222x0 \ALUSHT/SHT/U908  ( .ZN(\ALUSHT/SHT/n2738 ), .A(
        \ALUSHT/SHT/n3029 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n2403 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n3031 ), .F(\ALUSHT/SHT/n2454 )
         );
    snl_oai222x0 \ALUSHT/SHT/U1014  ( .ZN(\ALUSHT/SHT/n2486 ), .A(
        \ALUSHT/SHT/n2954 ), .B(\ALUSHT/SHT/n2402 ), .C(\ALUSHT/SHT/n2446 ), 
        .D(\ALUSHT/SHT/n2392 ), .E(\ALUSHT/SHT/n3036 ), .F(\ALUSHT/SHT/n2386 )
         );
    snl_invx05 \ALUSHT/SHT/U546  ( .ZN(\ALUSHT/SHT/n2520 ), .A(\pgaluina[4] )
         );
    snl_oa022x1 \ALUSHT/SHT/U561  ( .Z(\ALUSHT/SHT/n2543 ), .A(
        \ALUSHT/SHT/n2544 ), .B(\ALUSHT/SHT/n2502 ), .C(\ALUSHT/SHT/n2545 ), 
        .D(\ALUSHT/SHT/n2380 ) );
    snl_oai122x0 \ALUSHT/SHT/U883  ( .ZN(\ALUSHT/SHT/n2489 ), .A(
        \ALUSHT/SHT/n2516 ), .B(\ALUSHT/SHT/n2413 ), .C(\ALUSHT/SHT/n2961 ), 
        .D(\ALUSHT/SHT/n2382 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_oai2222x0 \ALUSHT/SHT/U913  ( .ZN(\ALUSHT/SHT/n2839 ), .A(
        \ALUSHT/SHT/n3011 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n3015 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3013 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3012 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_aoi222x0 \ALUSHT/SHT/U1028  ( .ZN(\ALUSHT/SHT/n3091 ), .A(
        \ALUSHT/SHT/n2421 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n3092 ), 
        .D(\ALUSHT/SHT/n2663 ), .E(\ALUSHT/SHT/n3063 ), .F(\ALUSHT/SHT/n2298 )
         );
    snl_aoi2222x1 \ALUSHT/SHT/U395  ( .ZN(\ALUSHT/SHT/n2921 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[15] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[16] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[17] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[14] ) );
    snl_aoi222x2 \ALUSHT/SHT/U433  ( .ZN(\ALUSHT/SHT/n2947 ), .A(
        \ALUSHT/SHT/n2946 ), .B(\ALUSHT/SHT/n2539 ), .C(\ALUSHT/SHT/n2778 ), 
        .D(\ALUSHT/SHT/n2694 ), .E(\ALUSHT/SHT/n2779 ), .F(\phshtd[2] ) );
    snl_aoi012x1 \ALUSHT/SHT/U676  ( .ZN(\ALUSHT/SHT/n2772 ), .A(
        \ALUSHT/SHT/n2423 ), .B(\pgaluina[23] ), .C(\ALUSHT/SHT/n2419 ) );
    snl_aoi122x0 \ALUSHT/SHT/U934  ( .ZN(\ALUSHT/SHT/n2691 ), .A(
        \ALUSHT/SHT/n2992 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n2988 ), 
        .D(\ALUSHT/SHT/n2298 ), .E(\ALUSHT/SHT/n2742 ) );
    snl_ao012x1 \ALUSHT/SHT/U808  ( .Z(\ALUSHT/SHT/n2949 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[11] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_oai122x0 \ALUSHT/SHT/U998  ( .ZN(\ALUSHT/SHT/n3076 ), .A(
        \ALUSHT/SHT/n3023 ), .B(\ALUSHT/SHT/n2657 ), .C(\ALUSHT/SHT/n3021 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n2764 ) );
    snl_oai222x0 \ALUSHT/SHT/U1084  ( .ZN(\ALUSHT/SHT/n2902 ), .A(
        \ALUSHT/SHT/n3080 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n2533 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n3094 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_invx05 \ALUSHT/SHT/U1114  ( .ZN(\ALUSHT/SHT/n3105 ), .A(
        \ALUSHT/SHT/n2979 ) );
    snl_oai122x0 \ALUSHT/SHT/U584  ( .ZN(\ALUSHT/SHT/n2604 ), .A(
        \ALUSHT/SHT/n2574 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2572 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi222x0 \ALUSHT/SHT/U693  ( .ZN(\ALUSHT/SHT/n2342 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2858 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2859 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2851 )
         );
    snl_nand02x1 \ALUSHT/SHT/U703  ( .ZN(\ALUSHT/SHT/n2415 ), .A(
        \ALUSHT/SHT/n2909 ), .B(\phshtd[5] ) );
    snl_oa222x1 \ALUSHT/SHT/U841  ( .Z(\ALUSHT/SHT/n2986 ), .A(
        \ALUSHT/SHT/n2985 ), .B(\ALUSHT/SHT/n2627 ), .C(\ALUSHT/SHT/n2984 ), 
        .D(\ALUSHT/SHT/n2638 ), .E(\ALUSHT/SHT/n2298 ), .F(\ALUSHT/SHT/n2983 )
         );
    snl_invx05 \ALUSHT/SHT/U724  ( .ZN(\ALUSHT/SHT/n2721 ), .A(
        \ALUSHT/SHT/n2621 ) );
    snl_aoi222x2 \ALUSHT/SHT/U414  ( .ZN(\ALUSHT/SHT/n2546 ), .A(
        \ALUSHT/SHT/n2547 ), .B(\ALUSHT/SHT/n2498 ), .C(\ALUSHT/SHT/n2548 ), 
        .D(\ALUSHT/SHT/n2542 ), .E(\ALUSHT/SHT/n2549 ), .F(\ALUSHT/SHT/n2503 )
         );
    snl_aoi022x1 \ALUSHT/SHT/U866  ( .ZN(\ALUSHT/SHT/n3006 ), .A(
        \pgaluina[30] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[29] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1046  ( .ZN(\ALUSHT/SHT/n2841 ), .A(
        \ALUSHT/SHT/n3099 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3088 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3095 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3097 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_nor03x1 \ALUSHT/SHT/U387  ( .ZN(\ALUSHT/SHT/n2645 ), .A(\poshtfnc[1] ), 
        .B(\poshtfnc[2] ), .C(\poshtfnc[0] ) );
    snl_invx1 \ALUSHT/SHT/U421  ( .ZN(\ALUSHT/SHT/n2500 ), .A(\phshtd[1] ) );
    snl_nand02x1 \ALUSHT/SHT/U528  ( .ZN(\ALUSHT/SHT/n2454 ), .A(
        \ALUSHT/SHT/n2503 ), .B(\ALUSHT/SHT/n2427 ) );
    snl_nand02x1 \ALUSHT/SHT/U618  ( .ZN(\ALUSHT/SHT/n2642 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n2503 ) );
    snl_oai222x0 \ALUSHT/SHT/U788  ( .ZN(\ALUSHT/SHT/n2853 ), .A(
        \ALUSHT/SHT/n2933 ), .B(\ALUSHT/SHT/n2615 ), .C(\ALUSHT/SHT/n2932 ), 
        .D(\ALUSHT/SHT/n2614 ), .E(\phshtd[2] ), .F(\ALUSHT/SHT/n2936 ) );
    snl_oai122x0 \ALUSHT/SHT/U853  ( .ZN(\ALUSHT/SHT/n2470 ), .A(
        \ALUSHT/SHT/n2515 ), .B(\ALUSHT/SHT/n2413 ), .C(\ALUSHT/SHT/n2998 ), 
        .D(\ALUSHT/SHT/n2382 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_oai2222x0 \ALUSHT/SHT/U948  ( .ZN(\ALUSHT/SHT/n2753 ), .A(
        \ALUSHT/SHT/n3038 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3047 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n2466 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3026 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_oa222x1 \ALUSHT/SHT/U1054  ( .Z(\ALUSHT/SHT/n2462 ), .A(
        \ALUSHT/SHT/n3046 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n2457 ), 
        .D(\ALUSHT/SHT/n2499 ), .E(\ALUSHT/SHT/n3055 ), .F(\ALUSHT/SHT/n2500 )
         );
    snl_nand02x1 \ALUSHT/SHT/U1061  ( .ZN(\ALUSHT/SHT/n2869 ), .A(
        \ALUSHT/SHT/n2867 ), .B(\ALUSHT/SHT/n2866 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1073  ( .ZN(\ALUSHT/SHT/n2889 ), .A(
        \ALUSHT/SHT/n3074 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3108 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n3109 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3071 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_aoi222x0 \ALUSHT/SHT/U681  ( .ZN(\ALUSHT/SHT/n2798 ), .A(
        \ALUSHT/SHT/n2656 ), .B(\ALUSHT/SHT/n2799 ), .C(\ALUSHT/SHT/n2800 ), 
        .D(\ALUSHT/SHT/n2441 ), .E(\ALUSHT/SHT/n2655 ), .F(\ALUSHT/SHT/n2801 )
         );
    snl_invx05 \ALUSHT/SHT/U711  ( .ZN(\ALUSHT/SHT/n2468 ), .A(
        \ALUSHT/SHT/n2640 ) );
    snl_invx05 \ALUSHT/SHT/U736  ( .ZN(\ALUSHT/SHT/n2480 ), .A(
        \ALUSHT/SHT/n2455 ) );
    snl_aoi022x1 \ALUSHT/SHT/U874  ( .ZN(\ALUSHT/SHT/n3013 ), .A(
        \pgaluina[18] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[17] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_nand02x3 \ALUSHT/SHT/U406  ( .ZN(\ALUSHT/SHT/n2380 ), .A(
        \ALUSHT/SHT/n2382 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_nor02x1 \ALUSHT/SHT/U596  ( .ZN(\ALUSHT/SHT/n2495 ), .A(
        \ALUSHT/SHT/n2499 ), .B(\ALUSHT/SHT/n2620 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U758  ( .ZN(\ALUSHT/SHT/n2926 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[29] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[30] ), .E(\pgaluina[31] ), .F(\ALUSHT/SHT/n2506 ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[28] ) );
    snl_aoi022x1 \ALUSHT/SHT/U282  ( .ZN(\ALUSHT/SHT/n2774 ), .A(
        \ALUSHT/SHT/n2404 ), .B(\ALUSHT/SHT/n2775 ), .C(\ALUSHT/SHT/n2776 ), 
        .D(\ALUSHT/SHT/n2386 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U285  ( .ZN(\ALUSHT/SHT/n2525 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[7] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[8] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[9] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[6] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U287  ( .ZN(\ALUSHT/SHT/n2529 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[6] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[7] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[8] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[5] ) );
    snl_aoi012x1 \ALUSHT/SHT/U317  ( .ZN(\ALUSHT/SHT/n2490 ), .A(\pgaluina[0] 
        ), .B(\ALUSHT/SHT/n2491 ), .C(\ALUSHT/SHT/n2492 ) );
    snl_aoi122x0 \ALUSHT/SHT/U345  ( .ZN(\ALUSHT/SHT/n2335 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[8] ), .C(\pgaluina[16] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U362  ( .ZN(\ALUSHT/SHT/n2305 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2796 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2854 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[25] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[1] ) );
    snl_nand02x1 \ALUSHT/SHT/U468  ( .ZN(\ALUSHT/pkshtout[2] ), .A(
        \ALUSHT/SHT/n2307 ), .B(\ALUSHT/SHT/n2308 ) );
    snl_oa222x1 \ALUSHT/SHT/U573  ( .Z(\ALUSHT/SHT/n2586 ), .A(
        \ALUSHT/SHT/n2587 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2527 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2588 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_oai022x1 \ALUSHT/SHT/U643  ( .ZN(\ALUSHT/SHT/n2675 ), .A(
        \ALUSHT/SHT/n2676 ), .B(\ALUSHT/SHT/n2619 ), .C(\ALUSHT/SHT/n2425 ), 
        .D(\ALUSHT/SHT/n2615 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1096  ( .ZN(\ALUSHT/SHT/n2784 ), .A(
        \ALUSHT/SHT/n2593 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n3077 ), 
        .D(\phshtd[4] ) );
    snl_invx05 \ALUSHT/SHT/U1106  ( .ZN(\ALUSHT/SHT/n3107 ), .A(
        \ALUSHT/SHT/n2999 ) );
    snl_invx05 \ALUSHT/SHT/U1121  ( .ZN(\ALUSHT/SHT/n3048 ), .A(
        \ALUSHT/SHT/n3046 ) );
    snl_invx05 \ALUSHT/SHT/U891  ( .ZN(\ALUSHT/SHT/n3021 ), .A(
        \ALUSHT/SHT/n2877 ) );
    snl_oai2222x0 \ALUSHT/SHT/U901  ( .ZN(\ALUSHT/SHT/n2783 ), .A(
        \ALUSHT/SHT/n2648 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2671 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2649 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2647 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai2222x0 \ALUSHT/SHT/U926  ( .ZN(\ALUSHT/SHT/n2887 ), .A(
        \ALUSHT/SHT/n2932 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2939 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2938 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2933 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_invx1 \ALUSHT/SHT/U379  ( .ZN(\ALUSHT/SHT/n2661 ), .A(
        \ALUSHT/SHT/n2499 ) );
    snl_oai022x1 \ALUSHT/SHT/U554  ( .ZN(\ALUSHT/SHT/n2530 ), .A(
        \ALUSHT/SHT/n2531 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2532 ), 
        .D(\ALUSHT/SHT/n2399 ) );
    snl_oa222x1 \ALUSHT/SHT/U568  ( .Z(\ALUSHT/SHT/n2571 ), .A(
        \ALUSHT/SHT/n2572 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2573 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2574 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_and34x0 \ALUSHT/SHT/U664  ( .Z(\ALUSHT/SHT/n2718 ), .A(
        \ALUSHT/SHT/n2578 ), .B(\ALUSHT/SHT/n2575 ), .C(\ALUSHT/SHT/n2571 ), 
        .D(\ALUSHT/SHT/n2567 ) );
    snl_oai222x0 \ALUSHT/SHT/U1021  ( .ZN(\ALUSHT/SHT/n2803 ), .A(
        \ALUSHT/SHT/n3086 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2678 ), 
        .D(\ALUSHT/SHT/n2614 ), .E(\ALUSHT/SHT/n2679 ), .F(\ALUSHT/SHT/n2500 )
         );
    snl_aoi222x1 \ALUSHT/SHT/U454  ( .ZN(\ALUSHT/SHT/n2855 ), .A(
        \ALUSHT/SHT/n2662 ), .B(\ALUSHT/SHT/n2758 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2811 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2812 )
         );
    snl_nand04x0 \ALUSHT/SHT/U658  ( .ZN(\ALUSHT/SHT/n2712 ), .A(
        \ALUSHT/SHT/n2607 ), .B(\ALUSHT/SHT/n2608 ), .C(\ALUSHT/SHT/n2609 ), 
        .D(\ALUSHT/SHT/n2610 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U1006  ( .ZN(\ALUSHT/SHT/n3080 ), .A(
        \ALUSHT/SHT/n2386 ), .B(\ALUSHT/SHT/n2405 ), .C(\ALUSHT/SHT/n2658 ) );
    snl_oa2222x1 \ALUSHT/SHT/U764  ( .Z(\ALUSHT/SHT/n2582 ), .A(
        \ALUSHT/SHT/n2918 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2919 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2524 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2920 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_oai012x1 \ALUSHT/SHT/U826  ( .ZN(\ALUSHT/SHT/n2967 ), .A(
        \ALUSHT/SHT/n2518 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_nand02x1 \ALUSHT/SHT/U473  ( .ZN(\ALUSHT/pkshtout[7] ), .A(
        \ALUSHT/SHT/n2317 ), .B(\ALUSHT/SHT/n2318 ) );
    snl_ao122x1 \ALUSHT/SHT/U801  ( .Z(\ALUSHT/SHT/n2779 ), .A(\pgaluina[8] ), 
        .B(\ALUSHT/SHT/n2432 ), .C(\ALUSHT/SHT/n2427 ), .D(\ALUSHT/SHT/n2945 ), 
        .E(\ALUSHT/SHT/n2433 ) );
    snl_ao122x1 \ALUSHT/SHT/U991  ( .Z(\ALUSHT/SHT/n3072 ), .A(\pgaluina[9] ), 
        .B(\ALUSHT/SHT/n2432 ), .C(\ALUSHT/SHT/n2427 ), .D(\ALUSHT/SHT/n2956 ), 
        .E(\ALUSHT/SHT/n2433 ) );
    snl_invx05 \ALUSHT/SHT/U743  ( .ZN(\ALUSHT/SHT/n2389 ), .A(
        \ALUSHT/SHT/n2664 ) );
    snl_oai122x0 \ALUSHT/SHT/U848  ( .ZN(\ALUSHT/SHT/n2994 ), .A(
        \ALUSHT/SHT/n2513 ), .B(\ALUSHT/SHT/n2413 ), .C(\ALUSHT/SHT/n2993 ), 
        .D(\ALUSHT/SHT/n2382 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_oai122x0 \ALUSHT/SHT/U974  ( .ZN(\ALUSHT/SHT/n3065 ), .A(
        \ALUSHT/SHT/n2984 ), .B(\ALUSHT/SHT/n2627 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n3064 ), .E(\ALUSHT/SHT/n2772 ) );
    snl_nand02x1 \ALUSHT/SHT/U496  ( .ZN(\ALUSHT/pkshtout[30] ), .A(
        \ALUSHT/SHT/n2363 ), .B(\ALUSHT/SHT/n2364 ) );
    snl_nand02x2 \ALUSHT/SHT/U297  ( .ZN(\ALUSHT/SHT/n2388 ), .A(\phshtd[2] ), 
        .B(\ALUSHT/SHT/n2298 ) );
    snl_aoi223x0 \ALUSHT/SHT/U320  ( .ZN(\ALUSHT/SHT/n2434 ), .A(
        \ALUSHT/SHT/n2435 ), .B(\ALUSHT/SHT/n2436 ), .C(\ALUSHT/SHT/n2437 ), 
        .D(\ALUSHT/SHT/n2438 ), .E(\ALUSHT/SHT/n2439 ), .F(\ALUSHT/SHT/n2440 ), 
        .G(\ALUSHT/SHT/n2441 ) );
    snl_oa2222x1 \ALUSHT/SHT/U330  ( .Z(\ALUSHT/SHT/n2955 ), .A(
        \ALUSHT/SHT/n2954 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2953 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2951 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2952 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi012x1 \ALUSHT/SHT/U506  ( .ZN(\ALUSHT/SHT/n2403 ), .A(
        \ALUSHT/SHT/n2404 ), .B(\ALUSHT/SHT/n2405 ), .C(\ALUSHT/SHT/n2391 ) );
    snl_aoi222x0 \ALUSHT/SHT/U521  ( .ZN(\ALUSHT/SHT/n2482 ), .A(
        \ALUSHT/SHT/n2478 ), .B(\ALUSHT/SHT/n2483 ), .C(\ALUSHT/SHT/n2484 ), 
        .D(\ALUSHT/SHT/n2441 ), .E(\ALUSHT/SHT/n2485 ), .F(\ALUSHT/SHT/n2486 )
         );
    snl_and02x1 \ALUSHT/SHT/U611  ( .Z(\ALUSHT/SHT/n2635 ), .A(
        \ALUSHT/SHT/n2624 ), .B(\ALUSHT/SHT/n2381 ) );
    snl_nor02x1 \ALUSHT/SHT/U636  ( .ZN(\ALUSHT/SHT/n2660 ), .A(
        \ALUSHT/SHT/n2621 ), .B(\phshtd[5] ) );
    snl_oai122x0 \ALUSHT/SHT/U1068  ( .ZN(\ALUSHT/SHT/n2885 ), .A(
        \ALUSHT/SHT/n3029 ), .B(\ALUSHT/SHT/n2536 ), .C(\ALUSHT/SHT/n3077 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2880 ) );
    snl_oai012x1 \ALUSHT/SHT/U781  ( .ZN(\ALUSHT/SHT/n2407 ), .A(
        \ALUSHT/SHT/n2654 ), .B(\ALUSHT/SHT/n2500 ), .C(\ALUSHT/SHT/n2551 ) );
    snl_oai022x1 \ALUSHT/SHT/U953  ( .ZN(\ALUSHT/SHT/n2811 ), .A(
        \ALUSHT/SHT/n2668 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2620 ), 
        .D(\ALUSHT/SHT/n2619 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U355  ( .ZN(\ALUSHT/SHT/n2313 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2740 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2746 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[29] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[5] ) );
    snl_aoi022x4 \ALUSHT/SHT/U397  ( .ZN(\ALUSHT/SHT/n2648 ), .A(
        \pgaluina[14] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[13] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_oai122x0 \ALUSHT/SHT/U586  ( .ZN(\ALUSHT/SHT/n2606 ), .A(
        \ALUSHT/SHT/n2580 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2579 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_invx05 \ALUSHT/SHT/U726  ( .ZN(\ALUSHT/SHT/n2485 ), .A(
        \ALUSHT/SHT/n2630 ) );
    snl_oai2222x0 \ALUSHT/SHT/U958  ( .ZN(\ALUSHT/SHT/n2759 ), .A(
        \ALUSHT/SHT/n2933 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2940 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2939 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2938 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1063  ( .ZN(\ALUSHT/SHT/n2870 ), .A(
        \ALUSHT/SHT/n3106 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3098 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3100 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3103 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai122x0 \ALUSHT/SHT/U1044  ( .ZN(\ALUSHT/SHT/n2840 ), .A(
        \ALUSHT/SHT/n2570 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3034 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2838 ) );
    snl_oai222x0 \ALUSHT/SHT/U864  ( .ZN(\ALUSHT/SHT/n2728 ), .A(
        \ALUSHT/SHT/n3004 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n2535 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2496 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_aoi2222x2 \ALUSHT/SHT/U416  ( .ZN(\ALUSHT/SHT/n2324 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2902 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2903 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[2] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2726 ) );
    snl_aoi012x4 \ALUSHT/SHT/U431  ( .ZN(\ALUSHT/SHT/n2701 ), .A(
        \ALUSHT/SHT/n2694 ), .B(\ALUSHT/SHT/n2702 ), .C(\ALUSHT/SHT/n2696 ) );
    snl_oai122x0 \ALUSHT/SHT/U843  ( .ZN(\ALUSHT/SHT/n2988 ), .A(
        \ALUSHT/SHT/n2511 ), .B(\ALUSHT/SHT/n2413 ), .C(\ALUSHT/SHT/n2987 ), 
        .D(\ALUSHT/SHT/n2382 ), .E(\ALUSHT/SHT/n2415 ) );
    snl_nand02x1 \ALUSHT/SHT/U478  ( .ZN(\ALUSHT/pkshtout[12] ), .A(
        \ALUSHT/SHT/n2327 ), .B(\ALUSHT/SHT/n2328 ) );
    snl_aoi222x0 \ALUSHT/SHT/U691  ( .ZN(\ALUSHT/SHT/n2344 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2850 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2851 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2845 )
         );
    snl_invx05 \ALUSHT/SHT/U701  ( .ZN(\ALUSHT/SHT/n2376 ), .A(
        \ALUSHT/SHT/n2445 ) );
    snl_invx05 \ALUSHT/SHT/U748  ( .ZN(\ALUSHT/SHT/n2592 ), .A(
        \ALUSHT/SHT/n2473 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1086  ( .ZN(\ALUSHT/SHT/n2903 ), .A(
        \ALUSHT/SHT/n2947 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n2950 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n2955 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3109 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_invx05 \ALUSHT/SHT/U1116  ( .ZN(\ALUSHT/SHT/n2997 ), .A(
        \ALUSHT/SHT/n2412 ) );
    snl_invx05 \ALUSHT/SHT/U544  ( .ZN(\ALUSHT/SHT/n2518 ), .A(\pgaluina[6] )
         );
    snl_oai2222x0 \ALUSHT/SHT/U936  ( .ZN(\ALUSHT/SHT/n2804 ), .A(
        \ALUSHT/SHT/n2647 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2674 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2671 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2649 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_invx2 \ALUSHT/SHT/U369  ( .ZN(\ALUSHT/SHT/n2298 ), .A(
        \ALUSHT/SHT/n2427 ) );
    snl_nand02x2 \ALUSHT/SHT/U372  ( .ZN(\ALUSHT/SHT/n2619 ), .A(\phshtd[1] ), 
        .B(\ALUSHT/SHT/n2386 ) );
    snl_nor04x0 \ALUSHT/SHT/U653  ( .ZN(\ALUSHT/SHT/n2707 ), .A(
        \ALUSHT/SHT/n2703 ), .B(\ALUSHT/SHT/n2704 ), .C(\ALUSHT/SHT/n2705 ), 
        .D(\ALUSHT/SHT/n2706 ) );
    snl_oai022x1 \ALUSHT/SHT/U674  ( .ZN(\ALUSHT/SHT/n2424 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n2769 ), .C(\ALUSHT/SHT/n2770 ), 
        .D(\ALUSHT/SHT/n2627 ) );
    snl_ao012x1 \ALUSHT/SHT/U881  ( .Z(\ALUSHT/SHT/n2685 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[8] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_oai012x1 \ALUSHT/SHT/U911  ( .ZN(\ALUSHT/SHT/n3033 ), .A(
        \ALUSHT/SHT/n3005 ), .B(\ALUSHT/SHT/n2500 ), .C(\ALUSHT/SHT/n2540 ) );
    snl_oai222x0 \ALUSHT/SHT/U563  ( .ZN(\ALUSHT/SHT/n2553 ), .A(
        \ALUSHT/SHT/n2554 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2540 ), 
        .D(\ALUSHT/SHT/n2538 ), .E(\ALUSHT/SHT/n2555 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U1016  ( .ZN(\ALUSHT/SHT/n2795 ), .A(
        \ALUSHT/SHT/n2466 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3055 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n2464 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3047 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_invx1 \ALUSHT/SHT/U444  ( .ZN(\ALUSHT/SHT/n2386 ), .A(\phshtd[2] ) );
    snl_invx1 \ALUSHT/SHT/U463  ( .ZN(\ALUSHT/SHT/n2631 ), .A(
        \ALUSHT/SHT/n2508 ) );
    snl_oai012x1 \ALUSHT/SHT/U578  ( .ZN(\ALUSHT/SHT/n2598 ), .A(
        \ALUSHT/SHT/n2552 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2396 ) );
    snl_oai222x0 \ALUSHT/SHT/U648  ( .ZN(\ALUSHT/SHT/n2690 ), .A(
        \ALUSHT/SHT/n2691 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n2467 ), 
        .D(\ALUSHT/SHT/n2499 ), .E(\ALUSHT/SHT/n2692 ), .F(\ALUSHT/SHT/n2500 )
         );
    snl_oa012x1 \ALUSHT/SHT/U811  ( .Z(\ALUSHT/SHT/n2952 ), .A(
        \ALUSHT/SHT/n2449 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_invx05 \ALUSHT/SHT/U1031  ( .ZN(\ALUSHT/SHT/n3094 ), .A(
        \ALUSHT/SHT/n2818 ) );
    snl_oa012x1 \ALUSHT/SHT/U981  ( .Z(\ALUSHT/SHT/n3068 ), .A(
        \ALUSHT/SHT/n2514 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_oai2222x0 \ALUSHT/SHT/U753  ( .ZN(\ALUSHT/SHT/n2590 ), .A(
        \ALUSHT/SHT/n2398 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2401 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2921 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2400 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_oai2222x0 \ALUSHT/SHT/U774  ( .ZN(\ALUSHT/SHT/n2863 ), .A(
        \ALUSHT/SHT/n2920 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2524 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2393 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2523 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_aoi222x0 \ALUSHT/SHT/U836  ( .ZN(\ALUSHT/SHT/n2980 ), .A(
        \ALUSHT/SHT/n2981 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2979 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2978 )
         );
    snl_nand02x1 \ALUSHT/SHT/U601  ( .ZN(\ALUSHT/SHT/n2626 ), .A(
        \pgaluina[15] ), .B(\ALUSHT/SHT/n2372 ) );
    snl_aoi022x1 \ALUSHT/SHT/U791  ( .ZN(\ALUSHT/SHT/n2939 ), .A(
        \pgaluina[23] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[22] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_oai2222x0 \ALUSHT/SHT/U858  ( .ZN(\ALUSHT/SHT/n2725 ), .A(
        \ALUSHT/SHT/n3001 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2986 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2991 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2996 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai2222x0 \ALUSHT/SHT/U943  ( .ZN(\ALUSHT/SHT/n2751 ), .A(
        \ALUSHT/SHT/n3007 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3011 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3010 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3008 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_nand02x1 \ALUSHT/SHT/U531  ( .ZN(\ALUSHT/SHT/n2374 ), .A(\poshtfnc[1] 
        ), .B(\poshtfnc[2] ) );
    snl_aoi122x0 \ALUSHT/SHT/U964  ( .ZN(\ALUSHT/SHT/n3057 ), .A(
        \pgaluina[16] ), .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(
        \ALUSHT/SHT/n2960 ), .E(\ALUSHT/SHT/n2419 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1078  ( .ZN(\ALUSHT/SHT/n2895 ), .A(
        \ALUSHT/SHT/n2976 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3104 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2963 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2969 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_aoi022x1 \ALUSHT/SHT/U307  ( .ZN(\ALUSHT/SHT/n2668 ), .A(\pgaluina[3] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[2] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_oai222x0 \ALUSHT/SHT/U516  ( .ZN(\ALUSHT/SHT/n2450 ), .A(
        \ALUSHT/SHT/n2451 ), .B(\ALUSHT/SHT/n2452 ), .C(\ALUSHT/SHT/n2453 ), 
        .D(\ALUSHT/SHT/n2454 ), .E(\ALUSHT/SHT/n2455 ), .F(\ALUSHT/SHT/n2456 )
         );
    snl_aoi022x1 \ALUSHT/SHT/U315  ( .ZN(\ALUSHT/SHT/n2673 ), .A(\pgaluina[4] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[3] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_aoi222x0 \ALUSHT/SHT/U332  ( .ZN(\ALUSHT/SHT/n3026 ), .A(
        \ALUSHT/SHT/n2949 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2775 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2386 ), .F(\ALUSHT/SHT/n3024 )
         );
    snl_nand02x1 \ALUSHT/SHT/U486  ( .ZN(\ALUSHT/pkshtout[20] ), .A(
        \ALUSHT/SHT/n2343 ), .B(\ALUSHT/SHT/n2344 ) );
    snl_aoi022x1 \ALUSHT/SHT/U523  ( .ZN(\ALUSHT/SHT/n2493 ), .A(
        \ALUSHT/SHT/n2494 ), .B(\ALUSHT/SHT/n2427 ), .C(\ALUSHT/SHT/n2495 ), 
        .D(\ALUSHT/SHT/n2298 ) );
    snl_nand02x1 \ALUSHT/SHT/U613  ( .ZN(\ALUSHT/SHT/n2637 ), .A(
        \pgaluina[31] ), .B(\ALUSHT/SHT/n2372 ) );
    snl_oa022x1 \ALUSHT/SHT/U626  ( .Z(\ALUSHT/SHT/n2653 ), .A(
        \ALUSHT/SHT/n2618 ), .B(\ALUSHT/SHT/n2300 ), .C(\ALUSHT/SHT/n2654 ), 
        .D(\ALUSHT/SHT/n2301 ) );
    snl_oai222x0 \ALUSHT/SHT/U783  ( .ZN(\ALUSHT/SHT/n2722 ), .A(
        \ALUSHT/SHT/n2456 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n2534 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2493 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U951  ( .ZN(\ALUSHT/SHT/n2812 ), .A(
        \ALUSHT/SHT/n2617 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2669 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2670 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2667 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nand02x1 \ALUSHT/SHT/U494  ( .ZN(\ALUSHT/pkshtout[28] ), .A(
        \ALUSHT/SHT/n2359 ), .B(\ALUSHT/SHT/n2360 ) );
    snl_aoi012x1 \ALUSHT/SHT/U299  ( .ZN(\ALUSHT/SHT/n2953 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[14] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_oai022x1 \ALUSHT/SHT/U329  ( .ZN(\ALUSHT/SHT/n2818 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n3079 ), .C(\ALUSHT/SHT/n3030 ), 
        .D(\ALUSHT/SHT/n2402 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U347  ( .ZN(\ALUSHT/SHT/n2329 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2884 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2891 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[21] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[13] ) );
    snl_aoi222x2 \ALUSHT/SHT/U438  ( .ZN(\ALUSHT/SHT/n3055 ), .A(
        \ALUSHT/SHT/n2949 ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2408 ), 
        .D(\ALUSHT/SHT/n2539 ), .E(\ALUSHT/SHT/n3024 ), .F(\phshtd[2] ) );
    snl_nor02x1 \ALUSHT/SHT/U504  ( .ZN(\ALUSHT/SHT/n2391 ), .A(
        \ALUSHT/SHT/n2392 ), .B(\ALUSHT/SHT/n2393 ) );
    snl_oa022x1 \ALUSHT/SHT/U634  ( .Z(\ALUSHT/SHT/n2658 ), .A(
        \ALUSHT/SHT/n2647 ), .B(\ALUSHT/SHT/n2300 ), .C(\ALUSHT/SHT/n2648 ), 
        .D(\ALUSHT/SHT/n2301 ) );
    snl_oai012x1 \ALUSHT/SHT/U976  ( .ZN(\ALUSHT/SHT/n2421 ), .A(
        \ALUSHT/SHT/n2513 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_aoi222x0 \ALUSHT/SHT/U698  ( .ZN(\ALUSHT/SHT/n2886 ), .A(
        \ALUSHT/SHT/n2849 ), .B(\ALUSHT/SHT/n2843 ), .C(\ALUSHT/SHT/n2810 ), 
        .D(\ALUSHT/SHT/n2801 ), .E(\ALUSHT/SHT/n2662 ), .F(\ALUSHT/SHT/n2887 )
         );
    snl_invx05 \ALUSHT/SHT/U708  ( .ZN(\ALUSHT/SHT/n2537 ), .A(
        \ALUSHT/SHT/n2510 ) );
    snl_aoi222x1 \ALUSHT/SHT/U456  ( .ZN(\ALUSHT/SHT/n2846 ), .A(
        \ALUSHT/SHT/n2662 ), .B(\ALUSHT/SHT/n2750 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2806 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2804 )
         );
    snl_nand02x1 \ALUSHT/SHT/U471  ( .ZN(\ALUSHT/pkshtout[5] ), .A(
        \ALUSHT/SHT/n2313 ), .B(\ALUSHT/SHT/n2314 ) );
    snl_nand02x1 \ALUSHT/SHT/U741  ( .ZN(\ALUSHT/SHT/n2917 ), .A(\pgaluina[0] 
        ), .B(\ALUSHT/SHT/n2504 ) );
    snl_nand02x1 \ALUSHT/SHT/U803  ( .ZN(\ALUSHT/SHT/n2409 ), .A(\phshtd[4] ), 
        .B(\ALUSHT/SHT/n2374 ) );
    snl_invx05 \ALUSHT/SHT/U993  ( .ZN(\ALUSHT/SHT/n3074 ), .A(
        \ALUSHT/SHT/n3073 ) );
    snl_oa122x1 \ALUSHT/SHT/U766  ( .Z(\ALUSHT/SHT/n2564 ), .A(
        \ALUSHT/SHT/n2401 ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2397 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2701 ) );
    snl_oa2222x1 \ALUSHT/SHT/U824  ( .Z(\ALUSHT/SHT/n2963 ), .A(
        \ALUSHT/SHT/n2964 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2961 ), 
        .D(\ALUSHT/SHT/n2627 ), .E(\ALUSHT/SHT/n2962 ), .F(\ALUSHT/SHT/n2501 ), 
        .G(\ALUSHT/SHT/n2959 ), .H(\ALUSHT/SHT/n2638 ) );
    snl_invx05 \ALUSHT/SHT/U888  ( .ZN(\ALUSHT/SHT/n3020 ), .A(
        \ALUSHT/SHT/n2767 ) );
    snl_oai122x0 \ALUSHT/SHT/U918  ( .ZN(\ALUSHT/SHT/n3039 ), .A(
        \ALUSHT/SHT/n2968 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2966 ), 
        .D(\ALUSHT/SHT/n2427 ), .E(\ALUSHT/SHT/n2737 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1004  ( .ZN(\ALUSHT/SHT/n2861 ), .A(
        \ALUSHT/SHT/n2649 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2673 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2674 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2671 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_aoi222x0 \ALUSHT/SHT/U1023  ( .ZN(\ALUSHT/SHT/n3088 ), .A(
        \ALUSHT/SHT/n2417 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n3089 ), 
        .D(\ALUSHT/SHT/n2663 ), .E(\ALUSHT/SHT/n3056 ), .F(\ALUSHT/SHT/n2298 )
         );
    snl_aoi2222x0 \ALUSHT/SHT/U360  ( .ZN(\ALUSHT/SHT/n2307 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2762 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2797 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[26] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[2] ) );
    snl_oa022x1 \ALUSHT/SHT/U556  ( .Z(\ALUSHT/SHT/n2534 ), .A(
        \ALUSHT/SHT/n2525 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2395 ), 
        .D(\ALUSHT/SHT/n2399 ) );
    snl_oa222x1 \ALUSHT/SHT/U571  ( .Z(\ALUSHT/SHT/n2581 ), .A(
        \ALUSHT/SHT/n2387 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2533 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2582 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U641  ( .ZN(\ALUSHT/SHT/n2494 ), .A(
        \ALUSHT/SHT/n2667 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2668 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2669 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n2670 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nor04x0 \ALUSHT/SHT/U666  ( .ZN(\ALUSHT/SHT/n2720 ), .A(
        \ALUSHT/SHT/n2719 ), .B(\ALUSHT/SHT/n2543 ), .C(\ALUSHT/SHT/n2550 ), 
        .D(\ALUSHT/SHT/n2546 ) );
    snl_invx05 \ALUSHT/SHT/U924  ( .ZN(\ALUSHT/SHT/n3042 ), .A(
        \ALUSHT/SHT/n2801 ) );
    snl_oai122x0 \ALUSHT/SHT/U1038  ( .ZN(\ALUSHT/SHT/n2832 ), .A(
        \ALUSHT/SHT/n2577 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3009 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2828 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U385  ( .ZN(\ALUSHT/SHT/n2327 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2890 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2896 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[20] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[12] ) );
    snl_invx05 \ALUSHT/SHT/U734  ( .ZN(\ALUSHT/SHT/n2569 ), .A(
        \ALUSHT/SHT/n2391 ) );
    snl_oai012x1 \ALUSHT/SHT/U818  ( .ZN(\ALUSHT/SHT/n2960 ), .A(
        \ALUSHT/SHT/n2522 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_oai2222x0 \ALUSHT/SHT/U893  ( .ZN(\ALUSHT/SHT/n2835 ), .A(
        \ALUSHT/SHT/n2939 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2943 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2941 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2940 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai023x0 \ALUSHT/SHT/U903  ( .ZN(\ALUSHT/SHT/n2792 ), .A(
        \ALUSHT/SHT/n2522 ), .B(\ALUSHT/SHT/n2374 ), .C(\ALUSHT/SHT/n2508 ), 
        .D(\phshtd[1] ), .E(\ALUSHT/SHT/n2672 ) );
    snl_invx05 \ALUSHT/SHT/U988  ( .ZN(\ALUSHT/SHT/n2788 ), .A(
        \ALUSHT/SHT/n2365 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1094  ( .ZN(\ALUSHT/SHT/n3070 ), .A(
        \ALUSHT/SHT/n2677 ), .B(\ALUSHT/SHT/n2504 ), .C(\ALUSHT/SHT/n2675 ), 
        .D(\phshtd[0] ) );
    snl_invx05 \ALUSHT/SHT/U1104  ( .ZN(\ALUSHT/SHT/n3110 ), .A(
        \ALUSHT/SHT/n2530 ) );
    snl_nand02x2 \ALUSHT/SHT/U404  ( .ZN(\ALUSHT/SHT/n2399 ), .A(\phshtd[2] ), 
        .B(\ALUSHT/SHT/n2427 ) );
    snl_aoi122x2 \ALUSHT/SHT/U423  ( .ZN(\ALUSHT/SHT/n2355 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[2] ), .C(\pgaluina[26] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_oa022x1 \ALUSHT/SHT/U594  ( .Z(\ALUSHT/SHT/n2616 ), .A(
        \ALUSHT/SHT/n2617 ), .B(\ALUSHT/SHT/n2300 ), .C(\ALUSHT/SHT/n2618 ), 
        .D(\ALUSHT/SHT/n2301 ) );
    snl_invx05 \ALUSHT/SHT/U876  ( .ZN(\ALUSHT/SHT/n3014 ), .A(
        \ALUSHT/SHT/n2829 ) );
    snl_invx05 \ALUSHT/SHT/U538  ( .ZN(\ALUSHT/SHT/n2512 ), .A(\pgaluina[12] )
         );
    snl_aoi222x0 \ALUSHT/SHT/U683  ( .ZN(\ALUSHT/SHT/n2360 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2807 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2808 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2803 )
         );
    snl_aoi222x0 \ALUSHT/SHT/U851  ( .ZN(\ALUSHT/SHT/n2996 ), .A(
        \ALUSHT/SHT/n2997 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2995 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2994 )
         );
    snl_nand02x1 \ALUSHT/SHT/U713  ( .ZN(\ALUSHT/SHT/n2594 ), .A(
        \pgaluina[31] ), .B(\ALUSHT/SHT/n2498 ) );
    snl_oai222x0 \ALUSHT/SHT/U1071  ( .ZN(\ALUSHT/SHT/n2882 ), .A(
        \ALUSHT/SHT/n3031 ), .B(\ALUSHT/SHT/n2638 ), .C(\phshtd[4] ), .D(
        \ALUSHT/SHT/n2472 ), .E(\ALUSHT/SHT/n3029 ), .F(\ALUSHT/SHT/n2640 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U382  ( .ZN(\ALUSHT/SHT/n2319 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2725 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2731 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[16] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[8] ) );
    snl_invx1 \ALUSHT/SHT/U403  ( .ZN(\ALUSHT/SHT/n2404 ), .A(
        \ALUSHT/SHT/n2399 ) );
    snl_aoi122x2 \ALUSHT/SHT/U424  ( .ZN(\ALUSHT/SHT/n2361 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[5] ), .C(\pgaluina[29] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_nand02x1 \ALUSHT/SHT/U608  ( .ZN(\ALUSHT/SHT/n2632 ), .A(
        \ALUSHT/SHT/n2624 ), .B(exetype1) );
    snl_aoi2222x0 \ALUSHT/SHT/U1056  ( .ZN(\ALUSHT/SHT/n3103 ), .A(
        \ALUSHT/SHT/n2995 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n3092 ), 
        .D(\ALUSHT/SHT/n2428 ), .E(\ALUSHT/SHT/n2997 ), .F(\ALUSHT/SHT/n2663 ), 
        .G(\ALUSHT/SHT/n2421 ), .H(\ALUSHT/SHT/n2911 ) );
    snl_aoi222x0 \ALUSHT/SHT/U684  ( .ZN(\ALUSHT/SHT/n2358 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2815 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2816 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2808 )
         );
    snl_invx05 \ALUSHT/SHT/U714  ( .ZN(\ALUSHT/SHT/n2909 ), .A(
        \ALUSHT/SHT/n2637 ) );
    snl_invx05 \ALUSHT/SHT/U798  ( .ZN(\ALUSHT/SHT/n2944 ), .A(
        \ALUSHT/SHT/n2825 ) );
    snl_invx05 \ALUSHT/SHT/U856  ( .ZN(\ALUSHT/SHT/n2469 ), .A(
        \ALUSHT/SHT/n3000 ) );
    snl_nand02x1 \ALUSHT/SHT/U593  ( .ZN(\ALUSHT/SHT/n2613 ), .A(
        \ALUSHT/SHT/n2477 ), .B(\ALUSHT/SHT/n2504 ) );
    snl_aoi022x1 \ALUSHT/SHT/U871  ( .ZN(\ALUSHT/SHT/n3010 ), .A(
        \pgaluina[24] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[23] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi122x0 \ALUSHT/SHT/U518  ( .ZN(\ALUSHT/SHT/n2467 ), .A(
        \ALUSHT/SHT/n2468 ), .B(\ALUSHT/SHT/n2469 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n2470 ), .E(\ALUSHT/SHT/n2471 ) );
    snl_nor03x0 \ALUSHT/SHT/U733  ( .ZN(\ALUSHT/SHT/n2378 ), .A(
        \ALUSHT/SHT/n2455 ), .B(\phshtd[0] ), .C(\ALUSHT/SHT/n2499 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U1051  ( .ZN(\ALUSHT/SHT/n3102 ), .A(
        \ALUSHT/SHT/n2974 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n3089 ), 
        .D(\ALUSHT/SHT/n2428 ), .E(\ALUSHT/SHT/n2975 ), .F(\ALUSHT/SHT/n2663 ), 
        .G(\ALUSHT/SHT/n2417 ), .H(\ALUSHT/SHT/n2911 ) );
    snl_oai122x0 \ALUSHT/SHT/U1076  ( .ZN(\ALUSHT/SHT/n2896 ), .A(
        \ALUSHT/SHT/n3049 ), .B(\ALUSHT/SHT/n2536 ), .C(\ALUSHT/SHT/n3087 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2892 ) );
    snl_aoi022x1 \ALUSHT/SHT/U309  ( .ZN(\ALUSHT/SHT/n2617 ), .A(
        \pgaluina[11] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[10] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_nand02x1 \ALUSHT/SHT/U488  ( .ZN(\ALUSHT/pkshtout[22] ), .A(
        \ALUSHT/SHT/n2347 ), .B(\ALUSHT/SHT/n2348 ) );
    snl_aoi122x0 \ALUSHT/SHT/U340  ( .ZN(\ALUSHT/SHT/n2345 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[13] ), .C(\pgaluina[21] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi222x0 \ALUSHT/SHT/U367  ( .ZN(\ALUSHT/SHT/n2969 ), .A(
        \ALUSHT/SHT/n2970 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2967 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2971 )
         );
    snl_nor02x1 \ALUSHT/SHT/U628  ( .ZN(\ALUSHT/SHT/n2655 ), .A(
        \ALUSHT/SHT/n2638 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_invx05 \ALUSHT/SHT/U894  ( .ZN(\ALUSHT/SHT/n3023 ), .A(
        \ALUSHT/SHT/n2835 ) );
    snl_aoi012x1 \ALUSHT/SHT/U1018  ( .ZN(\ALUSHT/SHT/n3085 ), .A(
        \ALUSHT/SHT/n2935 ), .B(\ALUSHT/SHT/n2390 ), .C(\ALUSHT/SHT/n2475 ) );
    snl_invx05 \ALUSHT/SHT/U904  ( .ZN(\ALUSHT/SHT/n3030 ), .A(
        \ALUSHT/SHT/n2792 ) );
    snl_oai222x0 \ALUSHT/SHT/U551  ( .ZN(\ALUSHT/SHT/n2473 ), .A(
        \ALUSHT/SHT/n2523 ), .B(\ALUSHT/SHT/n2399 ), .C(\ALUSHT/SHT/n2393 ), 
        .D(\ALUSHT/SHT/n2402 ), .E(\ALUSHT/SHT/n2524 ), .F(\ALUSHT/SHT/n2392 )
         );
    snl_oai122x0 \ALUSHT/SHT/U576  ( .ZN(\ALUSHT/SHT/n2595 ), .A(
        \ALUSHT/SHT/n2544 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2545 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi223x0 \ALUSHT/SHT/U646  ( .ZN(\ALUSHT/SHT/n2684 ), .A(
        \ALUSHT/SHT/n2661 ), .B(\ALUSHT/SHT/n2685 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n2686 ), .E(\ALUSHT/SHT/n2687 ), .F(\ALUSHT/SHT/n2459 ), 
        .G(\ALUSHT/SHT/n2542 ) );
    snl_nand04x0 \ALUSHT/SHT/U661  ( .ZN(\ALUSHT/SHT/n2715 ), .A(
        \ALUSHT/SHT/n2591 ), .B(\ALUSHT/SHT/n2595 ), .C(\ALUSHT/SHT/n2596 ), 
        .D(\ALUSHT/SHT/n2598 ) );
    snl_oai222x0 \ALUSHT/SHT/U923  ( .ZN(\ALUSHT/SHT/n2801 ), .A(
        \ALUSHT/SHT/n2620 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n2668 ), 
        .D(\ALUSHT/SHT/n2619 ), .E(\ALUSHT/SHT/n2669 ), .F(\ALUSHT/SHT/n2302 )
         );
    snl_aoi222x1 \ALUSHT/SHT/U451  ( .ZN(\ALUSHT/SHT/n2842 ), .A(
        \ALUSHT/SHT/n2548 ), .B(\ALUSHT/SHT/n2843 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2801 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2799 )
         );
    snl_invx05 \ALUSHT/SHT/U823  ( .ZN(\ALUSHT/SHT/n2488 ), .A(
        \ALUSHT/SHT/n2962 ) );
    snl_oai012x1 \ALUSHT/SHT/U838  ( .ZN(\ALUSHT/SHT/n2982 ), .A(
        \ALUSHT/SHT/n2652 ), .B(\ALUSHT/SHT/n2366 ), .C(\ALUSHT/SHT/n2637 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1093  ( .ZN(\ALUSHT/SHT/n2766 ), .A(
        \ALUSHT/SHT/n2545 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n2544 ), 
        .D(\phshtd[4] ) );
    snl_invx05 \ALUSHT/SHT/U1103  ( .ZN(\ALUSHT/SHT/n2611 ), .A(
        \ALUSHT/SHT/n2590 ) );
    snl_nand02x1 \ALUSHT/SHT/U476  ( .ZN(\ALUSHT/pkshtout[10] ), .A(
        \ALUSHT/SHT/n2323 ), .B(\ALUSHT/SHT/n2324 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U746  ( .ZN(\ALUSHT/SHT/n2919 ), .A(
        \pgaluina[20] ), .B(\ALUSHT/SHT/n2631 ), .C(\pgaluina[21] ), .D(
        \ALUSHT/SHT/n2541 ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[22] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[19] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U761  ( .ZN(\ALUSHT/SHT/n2928 ), .A(
        \pgaluina[21] ), .B(\ALUSHT/SHT/n2631 ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[22] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[23] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[20] ) );
    snl_ao012x1 \ALUSHT/SHT/U804  ( .Z(\ALUSHT/SHT/n2946 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[12] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_oai122x0 \ALUSHT/SHT/U1088  ( .ZN(\ALUSHT/SHT/n2908 ), .A(
        \ALUSHT/SHT/n2490 ), .B(\ALUSHT/SHT/n2377 ), .C(\ALUSHT/SHT/n3084 ), 
        .D(\ALUSHT/SHT/n2508 ), .E(\ALUSHT/SHT/n3111 ) );
    snl_invx05 \ALUSHT/SHT/U1118  ( .ZN(\ALUSHT/SHT/n2981 ), .A(
        \ALUSHT/SHT/n2448 ) );
    snl_aoi222x0 \ALUSHT/SHT/U994  ( .ZN(\ALUSHT/SHT/n3075 ), .A(
        \ALUSHT/SHT/n3072 ), .B(\ALUSHT/SHT/n2682 ), .C(\ALUSHT/SHT/n2430 ), 
        .D(\ALUSHT/SHT/n2435 ), .E(\ALUSHT/SHT/n2500 ), .F(\ALUSHT/SHT/n3073 )
         );
    snl_nand12x1 \ALUSHT/SHT/U503  ( .ZN(\ALUSHT/SHT/n2384 ), .A(
        \ALUSHT/SHT/n2385 ), .B(\ALUSHT/SHT/n2386 ) );
    snl_oai022x1 \ALUSHT/SHT/U633  ( .ZN(\ALUSHT/SHT/n2367 ), .A(
        \ALUSHT/SHT/n2434 ), .B(\ALUSHT/SHT/n2632 ), .C(\ALUSHT/SHT/n2442 ), 
        .D(\ALUSHT/SHT/n2381 ) );
    snl_oai223x0 \ALUSHT/SHT/U938  ( .ZN(\ALUSHT/SHT/n2806 ), .A(
        \ALUSHT/SHT/n2301 ), .B(\ALUSHT/SHT/n2522 ), .C(\ALUSHT/SHT/n2613 ), 
        .D(\ALUSHT/SHT/n2672 ), .E(\ALUSHT/SHT/n2619 ), .F(\ALUSHT/SHT/n2673 ), 
        .G(\ALUSHT/SHT/n2499 ) );
    snl_oai222x0 \ALUSHT/SHT/U1003  ( .ZN(\ALUSHT/SHT/n2787 ), .A(
        \ALUSHT/SHT/n3078 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2676 ), 
        .D(\ALUSHT/SHT/n2614 ), .E(\ALUSHT/SHT/n3060 ), .F(\ALUSHT/SHT/n2500 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U1024  ( .ZN(\ALUSHT/SHT/n2808 ), .A(
        \ALUSHT/SHT/n3088 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2676 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3059 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3078 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oa122x1 \ALUSHT/SHT/U971  ( .Z(\ALUSHT/SHT/n2678 ), .A(
        \ALUSHT/SHT/n3062 ), .B(\ALUSHT/SHT/n2627 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n3061 ), .E(\ALUSHT/SHT/n2771 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U290  ( .ZN(\ALUSHT/SHT/n2395 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[3] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[4] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[5] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[2] ) );
    snl_aoi012x1 \ALUSHT/SHT/U300  ( .ZN(\ALUSHT/SHT/n2446 ), .A(\pgaluina[2] 
        ), .B(\ALUSHT/SHT/n2409 ), .C(\ALUSHT/SHT/n2410 ) );
    snl_aoi223x0 \ALUSHT/SHT/U312  ( .ZN(\ALUSHT/SHT/n2476 ), .A(\pgaluina[0] 
        ), .B(\ALUSHT/SHT/n2477 ), .C(\ALUSHT/SHT/n2478 ), .D(
        \ALUSHT/SHT/n2437 ), .E(\ALUSHT/SHT/n2479 ), .F(\ALUSHT/SHT/n2480 ), 
        .G(\ALUSHT/SHT/n2481 ) );
    snl_nand02x1 \ALUSHT/SHT/U493  ( .ZN(\ALUSHT/pkshtout[27] ), .A(
        \ALUSHT/SHT/n2357 ), .B(\ALUSHT/SHT/n2358 ) );
    snl_aoi222x0 \ALUSHT/SHT/U335  ( .ZN(\ALUSHT/SHT/n3084 ), .A(
        \ALUSHT/SHT/n2978 ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2447 ), 
        .D(\ALUSHT/SHT/n2539 ), .E(\ALUSHT/SHT/n3039 ), .F(\phshtd[2] ) );
    snl_oai222x0 \ALUSHT/SHT/U956  ( .ZN(\ALUSHT/SHT/n2760 ), .A(
        \ALUSHT/SHT/n3052 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n3054 ), 
        .D(\ALUSHT/SHT/n2455 ), .E(\ALUSHT/SHT/n3053 ), .F(\ALUSHT/SHT/n2454 )
         );
    snl_aoi022x4 \ALUSHT/SHT/U399  ( .ZN(\ALUSHT/SHT/n2620 ), .A(\pgaluina[1] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[0] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_aoi2222x2 \ALUSHT/SHT/U418  ( .ZN(\ALUSHT/SHT/n2326 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2898 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2899 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[3] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2900 ) );
    snl_aoi022x1 \ALUSHT/SHT/U524  ( .ZN(\ALUSHT/SHT/n2496 ), .A(
        \ALUSHT/SHT/n2479 ), .B(\ALUSHT/SHT/n2427 ), .C(\ALUSHT/SHT/n2497 ), 
        .D(\ALUSHT/SHT/n2298 ) );
    snl_ao122x1 \ALUSHT/SHT/U588  ( .Z(\ALUSHT/SHT/n2608 ), .A(
        \ALUSHT/SHT/n2585 ), .B(\ALUSHT/SHT/n2537 ), .C(\ALUSHT/SHT/n2584 ), 
        .D(\ALUSHT/SHT/n2503 ), .E(\ALUSHT/SHT/n2597 ) );
    snl_nand02x1 \ALUSHT/SHT/U614  ( .ZN(\ALUSHT/SHT/n2638 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\phshtd[4] ) );
    snl_aoi022x1 \ALUSHT/SHT/U784  ( .ZN(\ALUSHT/SHT/n2932 ), .A(
        \pgaluina[29] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[28] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_nand02x1 \ALUSHT/SHT/U728  ( .ZN(\ALUSHT/SHT/n2913 ), .A(
        \ALUSHT/SHT/n2428 ), .B(\ALUSHT/SHT/n2483 ) );
    snl_nand02x1 \ALUSHT/SHT/U481  ( .ZN(\ALUSHT/pkshtout[15] ), .A(
        \ALUSHT/SHT/n2333 ), .B(\ALUSHT/SHT/n2334 ) );
    snl_oa222x1 \ALUSHT/SHT/U621  ( .Z(\ALUSHT/SHT/n2646 ), .A(
        \ALUSHT/SHT/n2647 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n2648 ), 
        .D(\ALUSHT/SHT/n2619 ), .E(\ALUSHT/SHT/n2649 ), .F(\ALUSHT/SHT/n2300 )
         );
    snl_oai012x1 \ALUSHT/SHT/U878  ( .ZN(\ALUSHT/SHT/n2831 ), .A(
        \ALUSHT/SHT/n3015 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2646 ) );
    snl_ao122x1 \ALUSHT/SHT/U511  ( .Z(\ALUSHT/SHT/n2420 ), .A(
        \ALUSHT/SHT/n2421 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n2418 ), 
        .D(\pgaluina[27] ), .E(\ALUSHT/SHT/n2419 ) );
    snl_oa2222x1 \ALUSHT/SHT/U327  ( .Z(\ALUSHT/SHT/n2544 ), .A(
        \ALUSHT/SHT/n2930 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2531 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2558 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2532 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_invx05 \ALUSHT/SHT/U536  ( .ZN(\ALUSHT/SHT/n2397 ), .A(\pgaluina[30] )
         );
    snl_ao122x1 \ALUSHT/SHT/U963  ( .Z(\ALUSHT/SHT/n3056 ), .A(\pgaluina[20] ), 
        .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(\ALUSHT/SHT/n2974 ), 
        .E(\ALUSHT/SHT/n2419 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U349  ( .ZN(\ALUSHT/SHT/n2321 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2726 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2727 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[17] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[9] ) );
    snl_nand02x1 \ALUSHT/SHT/U606  ( .ZN(\ALUSHT/SHT/n2463 ), .A(
        \ALUSHT/SHT/n2541 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_oai2222x0 \ALUSHT/SHT/U944  ( .ZN(\ALUSHT/SHT/n2749 ), .A(
        \ALUSHT/SHT/n3012 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2648 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3015 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3013 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_nand02x1 \ALUSHT/SHT/U1058  ( .ZN(\ALUSHT/SHT/n2864 ), .A(
        \ALUSHT/SHT/n2862 ), .B(\ALUSHT/SHT/n2860 ) );
    snl_aoi022x1 \ALUSHT/SHT/U796  ( .ZN(\ALUSHT/SHT/n2943 ), .A(
        \pgaluina[17] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[16] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi022x4 \ALUSHT/SHT/U443  ( .ZN(\ALUSHT/SHT/n2777 ), .A(
        \ALUSHT/SHT/n2404 ), .B(\ALUSHT/SHT/n2778 ), .C(\ALUSHT/SHT/n2779 ), 
        .D(\ALUSHT/SHT/n2386 ) );
    snl_nand02x1 \ALUSHT/SHT/U558  ( .ZN(\ALUSHT/SHT/n2536 ), .A(
        \ALUSHT/SHT/n2537 ), .B(\ALUSHT/SHT/n2427 ) );
    snl_ao012x1 \ALUSHT/SHT/U668  ( .Z(\ALUSHT/SHT/n2742 ), .A(
        \ALUSHT/SHT/n2651 ), .B(\pgaluina[5] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oa222x1 \ALUSHT/SHT/U1036  ( .Z(\ALUSHT/SHT/n3096 ), .A(
        \ALUSHT/SHT/n3062 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2998 ), 
        .D(\ALUSHT/SHT/n2501 ), .E(\ALUSHT/SHT/n3061 ), .F(\ALUSHT/SHT/n2427 )
         );
    snl_oai122x0 \ALUSHT/SHT/U1011  ( .ZN(\ALUSHT/SHT/n2819 ), .A(
        \ALUSHT/SHT/n3015 ), .B(\ALUSHT/SHT/n2619 ), .C(\ALUSHT/SHT/n3013 ), 
        .D(\ALUSHT/SHT/n2499 ), .E(\ALUSHT/SHT/n2658 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U754  ( .ZN(\ALUSHT/SHT/n2922 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[26] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[27] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[28] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[25] ) );
    snl_oa122x1 \ALUSHT/SHT/U773  ( .Z(\ALUSHT/SHT/n2554 ), .A(
        \ALUSHT/SHT/n2919 ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2664 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2693 ) );
    snl_ao012x1 \ALUSHT/SHT/U831  ( .Z(\ALUSHT/SHT/n2975 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[20] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U283  ( .ZN(\ALUSHT/SHT/n2531 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[9] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[10] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[11] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[8] ) );
    snl_aoi022x1 \ALUSHT/SHT/U313  ( .ZN(\ALUSHT/SHT/n2671 ), .A(\pgaluina[8] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[7] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_aoi2222x0 \ALUSHT/SHT/U352  ( .ZN(\ALUSHT/SHT/n2318 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2733 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2734 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[15] ), 
        .G(\ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2735 ) );
    snl_invx1 \ALUSHT/SHT/U375  ( .ZN(\ALUSHT/SHT/n2301 ), .A(
        \ALUSHT/SHT/n2686 ) );
    snl_aoi222x2 \ALUSHT/SHT/U458  ( .ZN(\ALUSHT/SHT/n2809 ), .A(
        \ALUSHT/SHT/n2810 ), .B(\ALUSHT/SHT/n2757 ), .C(\ALUSHT/SHT/n2655 ), 
        .D(\ALUSHT/SHT/n2811 ), .E(\ALUSHT/SHT/n2656 ), .F(\ALUSHT/SHT/n2812 )
         );
    snl_invx1 \ALUSHT/SHT/U464  ( .ZN(\ALUSHT/SHT/n2650 ), .A(
        \ALUSHT/SHT/n2613 ) );
    snl_oai2222x0 \ALUSHT/SHT/U768  ( .ZN(\ALUSHT/SHT/n2848 ), .A(
        \ALUSHT/SHT/n2924 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2925 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2529 ), .F(\ALUSHT/SHT/n2388 ), 
        .G(\ALUSHT/SHT/n2528 ), .H(\ALUSHT/SHT/n2402 ) );
    snl_oai2222x0 \ALUSHT/SHT/U816  ( .ZN(\ALUSHT/SHT/n2724 ), .A(
        \ALUSHT/SHT/n2950 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n2955 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n2958 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n2947 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_oai112x0 \ALUSHT/SHT/U986  ( .ZN(\ALUSHT/SHT/n2780 ), .A(
        \ALUSHT/SHT/n3060 ), .B(\ALUSHT/SHT/n2507 ), .C(\ALUSHT/SHT/n3069 ), 
        .D(\ALUSHT/SHT/n3070 ) );
    snl_oai122x0 \ALUSHT/SHT/U1081  ( .ZN(\ALUSHT/SHT/n2901 ), .A(
        \ALUSHT/SHT/n3052 ), .B(\ALUSHT/SHT/n2536 ), .C(\ALUSHT/SHT/n3090 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n2897 ) );
    snl_invx05 \ALUSHT/SHT/U1111  ( .ZN(\ALUSHT/SHT/n3037 ), .A(
        \ALUSHT/SHT/n2953 ) );
    snl_oai222x0 \ALUSHT/SHT/U564  ( .ZN(\ALUSHT/SHT/n2556 ), .A(
        \ALUSHT/SHT/n2557 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2558 ), 
        .D(\ALUSHT/SHT/n2538 ), .E(\ALUSHT/SHT/n2559 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_nor04x0 \ALUSHT/SHT/U654  ( .ZN(\ALUSHT/SHT/n2708 ), .A(
        \ALUSHT/SHT/n2595 ), .B(\ALUSHT/SHT/n2596 ), .C(\ALUSHT/SHT/n2598 ), 
        .D(\ALUSHT/SHT/n2599 ) );
    snl_invx05 \ALUSHT/SHT/U886  ( .ZN(\ALUSHT/SHT/n3019 ), .A(
        \ALUSHT/SHT/n2765 ) );
    snl_oa222x1 \ALUSHT/SHT/U916  ( .Z(\ALUSHT/SHT/n3038 ), .A(
        \ALUSHT/SHT/n2954 ), .B(\ALUSHT/SHT/n2399 ), .C(\ALUSHT/SHT/n2952 ), 
        .D(\ALUSHT/SHT/n2388 ), .E(\phshtd[2] ), .F(\ALUSHT/SHT/n3036 ) );
    snl_aoi012x1 \ALUSHT/SHT/U673  ( .ZN(\ALUSHT/SHT/n2768 ), .A(
        \ALUSHT/SHT/n2423 ), .B(\pgaluina[24] ), .C(\ALUSHT/SHT/n2419 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U390  ( .ZN(\ALUSHT/SHT/n2528 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[10] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[11] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[12] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[9] ) );
    snl_aoi222x1 \ALUSHT/SHT/U411  ( .ZN(\ALUSHT/SHT/n2867 ), .A(
        \ALUSHT/SHT/n2498 ), .B(\ALUSHT/SHT/n2868 ), .C(\ALUSHT/SHT/n2849 ), 
        .D(\ALUSHT/SHT/n2823 ), .E(\ALUSHT/SHT/n2548 ), .F(\ALUSHT/SHT/n2825 )
         );
    snl_aoi222x2 \ALUSHT/SHT/U436  ( .ZN(\ALUSHT/SHT/n3108 ), .A(
        \ALUSHT/SHT/n3037 ), .B(\ALUSHT/SHT/n2539 ), .C(\ALUSHT/SHT/n2681 ), 
        .D(\ALUSHT/SHT/n2694 ), .E(\ALUSHT/SHT/n2683 ), .F(\phshtd[2] ) );
    snl_invx05 \ALUSHT/SHT/U543  ( .ZN(\ALUSHT/SHT/n2517 ), .A(\pgaluina[7] )
         );
    snl_aoi222x0 \ALUSHT/SHT/U696  ( .ZN(\ALUSHT/SHT/n2336 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2874 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2875 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2870 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U931  ( .ZN(\ALUSHT/SHT/n2746 ), .A(
        \ALUSHT/SHT/n3044 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3042 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n3041 ), .F(\ALUSHT/SHT/n2642 ), 
        .G(\ALUSHT/SHT/n3045 ), .H(\ALUSHT/SHT/n2454 ) );
    snl_aoi122x0 \ALUSHT/SHT/U978  ( .ZN(\ALUSHT/SHT/n2769 ), .A(
        \pgaluina[21] ), .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(
        \ALUSHT/SHT/n2989 ), .E(\ALUSHT/SHT/n2419 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1043  ( .ZN(\ALUSHT/SHT/n2837 ), .A(
        \ALUSHT/SHT/n3098 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3086 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3091 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3096 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_nand02x1 \ALUSHT/SHT/U1064  ( .ZN(\ALUSHT/SHT/n2874 ), .A(
        \ALUSHT/SHT/n2873 ), .B(\ALUSHT/SHT/n2871 ) );
    snl_invx05 \ALUSHT/SHT/U706  ( .ZN(\ALUSHT/SHT/n2498 ), .A(
        \ALUSHT/SHT/n2380 ) );
    snl_oai012x1 \ALUSHT/SHT/U844  ( .ZN(\ALUSHT/SHT/n2989 ), .A(
        \ALUSHT/SHT/n2519 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_oai122x0 \ALUSHT/SHT/U581  ( .ZN(\ALUSHT/SHT/n2601 ), .A(
        \ALUSHT/SHT/n2562 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2561 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_nor02x1 \ALUSHT/SHT/U632  ( .ZN(\ALUSHT/SHT/n2423 ), .A(
        \ALUSHT/SHT/n2642 ), .B(\ALUSHT/SHT/n2374 ) );
    snl_invx05 \ALUSHT/SHT/U721  ( .ZN(\ALUSHT/SHT/n2810 ), .A(
        \ALUSHT/SHT/n2657 ) );
    snl_invx05 \ALUSHT/SHT/U863  ( .ZN(\ALUSHT/SHT/n3004 ), .A(
        \ALUSHT/SHT/n2481 ) );
    snl_oa012x1 \ALUSHT/SHT/U970  ( .Z(\ALUSHT/SHT/n3062 ), .A(
        \ALUSHT/SHT/n2515 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_nand02x1 \ALUSHT/SHT/U492  ( .ZN(\ALUSHT/pkshtout[26] ), .A(
        \ALUSHT/SHT/n2355 ), .B(\ALUSHT/SHT/n2356 ) );
    snl_aoi122x0 \ALUSHT/SHT/U298  ( .ZN(\ALUSHT/SHT/n3036 ), .A(\pgaluina[6] 
        ), .B(\ALUSHT/SHT/n2459 ), .C(\ALUSHT/SHT/n3037 ), .D(
        \ALUSHT/SHT/n2298 ), .E(\ALUSHT/SHT/n2460 ) );
    snl_aoi022x1 \ALUSHT/SHT/U308  ( .ZN(\ALUSHT/SHT/n2667 ), .A(\pgaluina[9] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[8] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_aoi222x0 \ALUSHT/SHT/U334  ( .ZN(\ALUSHT/SHT/n2852 ), .A(
        \ALUSHT/SHT/n2437 ), .B(\ALUSHT/SHT/n2823 ), .C(\ALUSHT/SHT/n2495 ), 
        .D(\ALUSHT/SHT/n2548 ), .E(\ALUSHT/SHT/n2480 ), .F(\ALUSHT/SHT/n2853 )
         );
    snl_nor02x1 \ALUSHT/SHT/U502  ( .ZN(\ALUSHT/SHT/n2383 ), .A(\phshtd[5] ), 
        .B(\ALUSHT/SHT/n2366 ) );
    snl_nand02x1 \ALUSHT/SHT/U525  ( .ZN(\ALUSHT/SHT/n2370 ), .A(\poshtfnc[2] 
        ), .B(\ALUSHT/SHT/n2372 ) );
    snl_oai222x0 \ALUSHT/SHT/U957  ( .ZN(\ALUSHT/SHT/n2758 ), .A(
        \ALUSHT/SHT/n2932 ), .B(\ALUSHT/SHT/n2615 ), .C(\ALUSHT/SHT/n2934 ), 
        .D(\ALUSHT/SHT/n2614 ), .E(\phshtd[2] ), .F(\ALUSHT/SHT/n2558 ) );
    snl_aoi122x0 \ALUSHT/SHT/U341  ( .ZN(\ALUSHT/SHT/n2343 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[12] ), .C(\pgaluina[20] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi222x0 \ALUSHT/SHT/U366  ( .ZN(\ALUSHT/SHT/n2976 ), .A(
        \ALUSHT/SHT/n2975 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2974 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2973 )
         );
    snl_aoi022x4 \ALUSHT/SHT/U398  ( .ZN(\ALUSHT/SHT/n2649 ), .A(
        \pgaluina[10] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[9] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_nand02x1 \ALUSHT/SHT/U615  ( .ZN(\ALUSHT/SHT/n2413 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\ALUSHT/SHT/n2382 ) );
    snl_invx05 \ALUSHT/SHT/U729  ( .ZN(\ALUSHT/SHT/n2433 ), .A(
        \ALUSHT/SHT/n2913 ) );
    snl_aoi022x1 \ALUSHT/SHT/U785  ( .ZN(\ALUSHT/SHT/n2933 ), .A(
        \pgaluina[27] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[26] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi2222x2 \ALUSHT/SHT/U419  ( .ZN(\ALUSHT/SHT/n2322 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2722 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2724 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[1] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2725 ) );
    snl_aoi222x1 \ALUSHT/SHT/U450  ( .ZN(\ALUSHT/SHT/n2866 ), .A(
        \ALUSHT/SHT/n2662 ), .B(\ALUSHT/SHT/n2853 ), .C(\ALUSHT/SHT/n2656 ), 
        .D(\ALUSHT/SHT/n2495 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2494 )
         );
    snl_oai122x0 \ALUSHT/SHT/U589  ( .ZN(\ALUSHT/SHT/n2609 ), .A(
        \ALUSHT/SHT/n2588 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2587 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi012x1 \ALUSHT/SHT/U822  ( .ZN(\ALUSHT/SHT/n2962 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[16] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_nand02x1 \ALUSHT/SHT/U477  ( .ZN(\ALUSHT/pkshtout[11] ), .A(
        \ALUSHT/SHT/n2325 ), .B(\ALUSHT/SHT/n2326 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U747  ( .ZN(\ALUSHT/SHT/n2920 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[16] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[17] ), .E(\pgaluina[18] ), .F(\ALUSHT/SHT/n2506 ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[15] ) );
    snl_invx05 \ALUSHT/SHT/U760  ( .ZN(\ALUSHT/SHT/n2698 ), .A(
        \ALUSHT/SHT/n2927 ) );
    snl_aoi012x1 \ALUSHT/SHT/U805  ( .ZN(\ALUSHT/SHT/n2948 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[15] ), .C(\ALUSHT/SHT/n2483 ) );
    snl_oai122x0 \ALUSHT/SHT/U995  ( .ZN(\ALUSHT/SHT/n2683 ), .A(
        \ALUSHT/SHT/n2514 ), .B(\ALUSHT/SHT/n2628 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n2952 ), .E(\ALUSHT/SHT/n2913 ) );
    snl_ao122x1 \ALUSHT/SHT/U577  ( .Z(\ALUSHT/SHT/n2596 ), .A(
        \ALUSHT/SHT/n2549 ), .B(\ALUSHT/SHT/n2537 ), .C(\ALUSHT/SHT/n2547 ), 
        .D(\ALUSHT/SHT/n2503 ), .E(\ALUSHT/SHT/n2597 ) );
    snl_oai2222x0 \ALUSHT/SHT/U895  ( .ZN(\ALUSHT/SHT/n2736 ), .A(
        \ALUSHT/SHT/n3022 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n3020 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n3019 ), .F(\ALUSHT/SHT/n2642 ), 
        .G(\ALUSHT/SHT/n3023 ), .H(\ALUSHT/SHT/n2454 ) );
    snl_oai222x0 \ALUSHT/SHT/U905  ( .ZN(\ALUSHT/SHT/n2785 ), .A(
        \ALUSHT/SHT/n2674 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2673 ), 
        .D(\ALUSHT/SHT/n2619 ), .E(\ALUSHT/SHT/n3030 ), .F(\ALUSHT/SHT/n2386 )
         );
    snl_invx05 \ALUSHT/SHT/U939  ( .ZN(\ALUSHT/SHT/n3050 ), .A(
        \ALUSHT/SHT/n2806 ) );
    snl_aoi012x1 \ALUSHT/SHT/U1025  ( .ZN(\ALUSHT/SHT/n3090 ), .A(
        \ALUSHT/SHT/n2758 ), .B(\ALUSHT/SHT/n2298 ), .C(\ALUSHT/SHT/n2530 ) );
    snl_nand04x0 \ALUSHT/SHT/U1089  ( .ZN(\ALUSHT/SHT/n2665 ), .A(
        \ALUSHT/SHT/n2709 ), .B(\ALUSHT/SHT/n2708 ), .C(\ALUSHT/SHT/n2711 ), 
        .D(\ALUSHT/SHT/n2707 ) );
    snl_invx05 \ALUSHT/SHT/U1119  ( .ZN(\ALUSHT/SHT/n2971 ), .A(
        \ALUSHT/SHT/n2966 ) );
    snl_aoi222x0 \ALUSHT/SHT/U1002  ( .ZN(\ALUSHT/SHT/n3078 ), .A(
        \ALUSHT/SHT/n2429 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n2965 ), 
        .D(\ALUSHT/SHT/n2663 ), .E(\ALUSHT/SHT/n2426 ), .F(\ALUSHT/SHT/n2298 )
         );
    snl_oai022x1 \ALUSHT/SHT/U647  ( .ZN(\ALUSHT/SHT/n2688 ), .A(
        \ALUSHT/SHT/n2689 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n2487 ), 
        .D(\ALUSHT/SHT/n2499 ) );
    snl_oai122x0 \ALUSHT/SHT/U1019  ( .ZN(\ALUSHT/SHT/n2802 ), .A(
        \ALUSHT/SHT/n3045 ), .B(\ALUSHT/SHT/n2657 ), .C(\ALUSHT/SHT/n3043 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n2798 ) );
    snl_nand04x0 \ALUSHT/SHT/U660  ( .ZN(\ALUSHT/SHT/n2714 ), .A(
        \ALUSHT/SHT/n2599 ), .B(\ALUSHT/SHT/n2600 ), .C(\ALUSHT/SHT/n2601 ), 
        .D(\ALUSHT/SHT/n2602 ) );
    snl_invx05 \ALUSHT/SHT/U922  ( .ZN(\ALUSHT/SHT/n3041 ), .A(
        \ALUSHT/SHT/n2799 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U383  ( .ZN(\ALUSHT/SHT/n2331 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2878 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2885 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[22] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[14] ) );
    snl_aoi122x2 \ALUSHT/SHT/U425  ( .ZN(\ALUSHT/SHT/n2351 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[0] ), .C(\pgaluina[24] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_invx05 \ALUSHT/SHT/U550  ( .ZN(\ALUSHT/SHT/n2522 ), .A(\pgaluina[0] )
         );
    snl_aoi222x0 \ALUSHT/SHT/U685  ( .ZN(\ALUSHT/SHT/n2356 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2820 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2821 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2816 )
         );
    snl_oa012x1 \ALUSHT/SHT/U839  ( .Z(\ALUSHT/SHT/n2984 ), .A(
        \ALUSHT/SHT/n2517 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_invx05 \ALUSHT/SHT/U1092  ( .ZN(\ALUSHT/SHT/n2830 ), .A(
        \ALUSHT/SHT/n2496 ) );
    snl_invx05 \ALUSHT/SHT/U1102  ( .ZN(\ALUSHT/SHT/n2584 ), .A(
        \ALUSHT/SHT/n2926 ) );
    snl_invx05 \ALUSHT/SHT/U715  ( .ZN(\ALUSHT/SHT/n2483 ), .A(
        \ALUSHT/SHT/n2626 ) );
    snl_aoi222x0 \ALUSHT/SHT/U857  ( .ZN(\ALUSHT/SHT/n3001 ), .A(
        \ALUSHT/SHT/n2469 ), .B(\ALUSHT/SHT/n2428 ), .C(\ALUSHT/SHT/n2999 ), 
        .D(\ALUSHT/SHT/n2911 ), .E(\ALUSHT/SHT/n2427 ), .F(\ALUSHT/SHT/n2470 )
         );
    snl_aoi0b12x0 \ALUSHT/SHT/U870  ( .ZN(\ALUSHT/SHT/n3009 ), .A(
        \ALUSHT/SHT/n2872 ), .B(\ALUSHT/SHT/n2298 ), .C(\ALUSHT/SHT/n2535 ) );
    snl_aoi2222x1 \ALUSHT/SHT/U402  ( .ZN(\ALUSHT/SHT/n2925 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[14] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[15] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[16] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[13] ) );
    snl_nand02x1 \ALUSHT/SHT/U592  ( .ZN(\ALUSHT/SHT/n2612 ), .A(\phshtd[0] ), 
        .B(\ALUSHT/SHT/n2477 ) );
    snl_nor02x1 \ALUSHT/SHT/U732  ( .ZN(\ALUSHT/SHT/n2696 ), .A(
        \ALUSHT/SHT/n2392 ), .B(\ALUSHT/SHT/n2366 ) );
    snl_nand02x1 \ALUSHT/SHT/U1050  ( .ZN(\ALUSHT/SHT/n2850 ), .A(
        \ALUSHT/SHT/n2847 ), .B(\ALUSHT/SHT/n2846 ) );
    snl_nand02x1 \ALUSHT/SHT/U489  ( .ZN(\ALUSHT/pkshtout[23] ), .A(
        \ALUSHT/SHT/n2349 ), .B(\ALUSHT/SHT/n2350 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U348  ( .ZN(\ALUSHT/SHT/n2323 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2900 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2904 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[18] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[10] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U353  ( .ZN(\ALUSHT/SHT/n2315 ), .A(
        \ALUSHT/SHT/n2641 ), .B(\ALUSHT/SHT/n2735 ), .C(\ALUSHT/SHT/n2643 ), 
        .D(\ALUSHT/SHT/n2741 ), .E(\ALUSHT/SHT/n2644 ), .F(\pgaluina[30] ), 
        .G(\ALUSHT/SHT/n2645 ), .H(\pgaluina[6] ) );
    snl_nand02x2 \ALUSHT/SHT/U374  ( .ZN(\ALUSHT/SHT/n2615 ), .A(\phshtd[2] ), 
        .B(\phshtd[1] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U391  ( .ZN(\ALUSHT/SHT/n2312 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2752 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2753 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[12] ), 
        .G(\ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2754 ) );
    snl_aoi122x2 \ALUSHT/SHT/U437  ( .ZN(\ALUSHT/SHT/n2579 ), .A(
        \pgaluina[30] ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2702 ), .D(
        \ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2914 ) );
    snl_aoi012x1 \ALUSHT/SHT/U519  ( .ZN(\ALUSHT/SHT/n2472 ), .A(
        \ALUSHT/SHT/n2390 ), .B(\ALUSHT/SHT/n2405 ), .C(\ALUSHT/SHT/n2473 ) );
    snl_nor02x1 \ALUSHT/SHT/U629  ( .ZN(\ALUSHT/SHT/n2656 ), .A(
        \ALUSHT/SHT/n2640 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1077  ( .ZN(\ALUSHT/SHT/n2894 ), .A(
        \ALUSHT/SHT/n3108 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3109 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n2947 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n3074 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_aoi222x0 \ALUSHT/SHT/U697  ( .ZN(\ALUSHT/SHT/n2880 ), .A(
        \ALUSHT/SHT/n2849 ), .B(\ALUSHT/SHT/n2839 ), .C(\ALUSHT/SHT/n2810 ), 
        .D(\ALUSHT/SHT/n2785 ), .E(\ALUSHT/SHT/n2662 ), .F(\ALUSHT/SHT/n2881 )
         );
    snl_invx05 \ALUSHT/SHT/U707  ( .ZN(\ALUSHT/SHT/n2435 ), .A(
        \ALUSHT/SHT/n2300 ) );
    snl_oa012x1 \ALUSHT/SHT/U979  ( .Z(\ALUSHT/SHT/n2770 ), .A(
        \ALUSHT/SHT/n2511 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_oa222x1 \ALUSHT/SHT/U1042  ( .Z(\ALUSHT/SHT/n3098 ), .A(
        \ALUSHT/SHT/n2984 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2985 ), 
        .D(\ALUSHT/SHT/n2501 ), .E(\ALUSHT/SHT/n3064 ), .F(\ALUSHT/SHT/n2427 )
         );
    snl_oai2222x0 \ALUSHT/SHT/U1065  ( .ZN(\ALUSHT/SHT/n2875 ), .A(
        \ALUSHT/SHT/n2963 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3099 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3102 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3104 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai122x0 \ALUSHT/SHT/U580  ( .ZN(\ALUSHT/SHT/n2600 ), .A(
        \ALUSHT/SHT/n2559 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2557 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi012x1 \ALUSHT/SHT/U845  ( .ZN(\ALUSHT/SHT/n2990 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[21] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_aoi222x1 \ALUSHT/SHT/U410  ( .ZN(\ALUSHT/SHT/n2847 ), .A(
        \ALUSHT/SHT/n2498 ), .B(\ALUSHT/SHT/n2848 ), .C(\ALUSHT/SHT/n2849 ), 
        .D(\ALUSHT/SHT/n2751 ), .E(\ALUSHT/SHT/n2548 ), .F(\ALUSHT/SHT/n2749 )
         );
    snl_aoi222x2 \ALUSHT/SHT/U459  ( .ZN(\ALUSHT/SHT/n2892 ), .A(
        \ALUSHT/SHT/n2849 ), .B(\ALUSHT/SHT/n2749 ), .C(\ALUSHT/SHT/n2810 ), 
        .D(\ALUSHT/SHT/n2806 ), .E(\ALUSHT/SHT/n2662 ), .F(\ALUSHT/SHT/n2751 )
         );
    snl_invx05 \ALUSHT/SHT/U720  ( .ZN(\ALUSHT/SHT/n2911 ), .A(
        \ALUSHT/SHT/n2638 ) );
    snl_oai012x1 \ALUSHT/SHT/U862  ( .ZN(\ALUSHT/SHT/n2481 ), .A(
        \ALUSHT/SHT/n3003 ), .B(\ALUSHT/SHT/n2499 ), .C(\ALUSHT/SHT/n2646 ) );
    snl_invx05 \ALUSHT/SHT/U769  ( .ZN(\ALUSHT/SHT/n2562 ), .A(
        \ALUSHT/SHT/n2848 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1080  ( .ZN(\ALUSHT/SHT/n2898 ), .A(
        \ALUSHT/SHT/n3053 ), .B(\ALUSHT/SHT/n2642 ), .C(\ALUSHT/SHT/n3052 ), 
        .D(\ALUSHT/SHT/n2454 ), .E(\ALUSHT/SHT/n3054 ), .F(\ALUSHT/SHT/n2451 ), 
        .G(\ALUSHT/SHT/n3110 ), .H(\ALUSHT/SHT/n2380 ) );
    snl_invx05 \ALUSHT/SHT/U1110  ( .ZN(\ALUSHT/SHT/n3081 ), .A(
        \ALUSHT/SHT/n3033 ) );
    snl_invx05 \ALUSHT/SHT/U542  ( .ZN(\ALUSHT/SHT/n2516 ), .A(\pgaluina[8] )
         );
    snl_oai222x0 \ALUSHT/SHT/U565  ( .ZN(\ALUSHT/SHT/n2560 ), .A(
        \ALUSHT/SHT/n2561 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2384 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n2562 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_nor04x0 \ALUSHT/SHT/U655  ( .ZN(\ALUSHT/SHT/n2709 ), .A(
        \ALUSHT/SHT/n2600 ), .B(\ALUSHT/SHT/n2601 ), .C(\ALUSHT/SHT/n2602 ), 
        .D(\ALUSHT/SHT/n2603 ) );
    snl_oai2222x0 \ALUSHT/SHT/U887  ( .ZN(\ALUSHT/SHT/n2767 ), .A(
        \ALUSHT/SHT/n2670 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2620 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2668 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2669 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_oai2222x0 \ALUSHT/SHT/U917  ( .ZN(\ALUSHT/SHT/n2739 ), .A(
        \ALUSHT/SHT/n3017 ), .B(\ALUSHT/SHT/n2630 ), .C(\ALUSHT/SHT/n3026 ), 
        .D(\ALUSHT/SHT/n2463 ), .E(\ALUSHT/SHT/n3038 ), .F(\ALUSHT/SHT/n2629 ), 
        .G(\ALUSHT/SHT/n2958 ), .H(\ALUSHT/SHT/n2465 ) );
    snl_aoi222x0 \ALUSHT/SHT/U672  ( .ZN(\ALUSHT/SHT/n2764 ), .A(
        \ALUSHT/SHT/n2656 ), .B(\ALUSHT/SHT/n2765 ), .C(\ALUSHT/SHT/n2766 ), 
        .D(\ALUSHT/SHT/n2441 ), .E(\ALUSHT/SHT/n2655 ), .F(\ALUSHT/SHT/n2767 )
         );
    snl_nand02x1 \ALUSHT/SHT/U559  ( .ZN(\ALUSHT/SHT/n2538 ), .A(
        \ALUSHT/SHT/n2537 ), .B(\ALUSHT/SHT/n2539 ) );
    snl_invx05 \ALUSHT/SHT/U930  ( .ZN(\ALUSHT/SHT/n3045 ), .A(
        \ALUSHT/SHT/n2843 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1037  ( .ZN(\ALUSHT/SHT/n2827 ), .A(
        \ALUSHT/SHT/n3096 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3066 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3086 ), .F(\ALUSHT/SHT/n2614 ), 
        .G(\ALUSHT/SHT/n3091 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_aoi2222x1 \ALUSHT/SHT/U442  ( .ZN(\ALUSHT/SHT/n2958 ), .A(
        \ALUSHT/SHT/n2458 ), .B(\ALUSHT/SHT/n2539 ), .C(\ALUSHT/SHT/n2957 ), 
        .D(\ALUSHT/SHT/n2404 ), .E(\ALUSHT/SHT/n2431 ), .F(\ALUSHT/SHT/n2390 ), 
        .G(\ALUSHT/SHT/n2956 ), .H(\ALUSHT/SHT/n2694 ) );
    snl_ao012x1 \ALUSHT/SHT/U669  ( .Z(\ALUSHT/SHT/n2747 ), .A(
        \ALUSHT/SHT/n2651 ), .B(\pgaluina[4] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_invx05 \ALUSHT/SHT/U1010  ( .ZN(\ALUSHT/SHT/n3082 ), .A(
        \ALUSHT/SHT/n2790 ) );
    snl_invx1 \ALUSHT/SHT/U465  ( .ZN(\ALUSHT/SHT/n2541 ), .A(
        \ALUSHT/SHT/n2507 ) );
    snl_invx05 \ALUSHT/SHT/U755  ( .ZN(\ALUSHT/SHT/n2700 ), .A(
        \ALUSHT/SHT/n2922 ) );
    snl_invx05 \ALUSHT/SHT/U772  ( .ZN(\ALUSHT/SHT/n2559 ), .A(
        \ALUSHT/SHT/n2857 ) );
    snl_oai012x1 \ALUSHT/SHT/U830  ( .ZN(\ALUSHT/SHT/n2974 ), .A(
        \ALUSHT/SHT/n2520 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U284  ( .ZN(\ALUSHT/SHT/n2523 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[8] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[9] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[10] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[7] ) );
    snl_aoi122x0 \ALUSHT/SHT/U291  ( .ZN(\ALUSHT/SHT/n2983 ), .A(
        \pgaluina[15] ), .B(\ALUSHT/SHT/n2915 ), .C(\ALUSHT/SHT/n2982 ), .D(
        \phshtd[4] ), .E(\ALUSHT/SHT/n2492 ) );
    snl_and02x1 \ALUSHT/SHT/U620  ( .Z(\ALUSHT/SHT/n2644 ), .A(
        \ALUSHT/SHT/n2633 ), .B(\ALUSHT/SHT/n2381 ) );
    snl_oa012x1 \ALUSHT/SHT/U817  ( .Z(\ALUSHT/SHT/n2959 ), .A(
        \ALUSHT/SHT/n2516 ), .B(\ALUSHT/SHT/n2636 ), .C(\ALUSHT/SHT/n2912 ) );
    snl_invx05 \ALUSHT/SHT/U879  ( .ZN(\ALUSHT/SHT/n3016 ), .A(
        \ALUSHT/SHT/n2831 ) );
    snl_nor02x1 \ALUSHT/SHT/U987  ( .ZN(\ALUSHT/SHT/n2365 ), .A(
        \ALUSHT/SHT/n2645 ), .B(\ALUSHT/SHT/n2634 ) );
    snl_aoi022x1 \ALUSHT/SHT/U296  ( .ZN(\ALUSHT/SHT/n2540 ), .A(
        \ALUSHT/SHT/n2541 ), .B(\pgaluina[1] ), .C(\ALUSHT/SHT/n2506 ), .D(
        \pgaluina[2] ) );
    snl_aoi012x1 \ALUSHT/SHT/U301  ( .ZN(\ALUSHT/SHT/n2954 ), .A(
        \ALUSHT/SHT/n2409 ), .B(\pgaluina[10] ), .C(\ALUSHT/SHT/n2410 ) );
    snl_ao122x1 \ALUSHT/SHT/U510  ( .Z(\ALUSHT/SHT/n2416 ), .A(
        \ALUSHT/SHT/n2417 ), .B(\ALUSHT/SHT/n2382 ), .C(\ALUSHT/SHT/n2418 ), 
        .D(\pgaluina[28] ), .E(\ALUSHT/SHT/n2419 ) );
    snl_aoi022x1 \ALUSHT/SHT/U306  ( .ZN(\ALUSHT/SHT/n2669 ), .A(\pgaluina[5] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[4] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_ao122x1 \ALUSHT/SHT/U321  ( .Z(\ALUSHT/SHT/n2807 ), .A(
        \ALUSHT/SHT/n2749 ), .B(\ALUSHT/SHT/n2810 ), .C(\ALUSHT/SHT/n2751 ), 
        .D(\ALUSHT/SHT/n2548 ), .E(\ALUSHT/SHT/n2297 ) );
    snl_aoi222x0 \ALUSHT/SHT/U326  ( .ZN(\ALUSHT/SHT/n2873 ), .A(
        \ALUSHT/SHT/n2498 ), .B(\ALUSHT/SHT/n2549 ), .C(\ALUSHT/SHT/n2849 ), 
        .D(\ALUSHT/SHT/n2829 ), .E(\ALUSHT/SHT/n2548 ), .F(\ALUSHT/SHT/n2831 )
         );
    snl_nand02x1 \ALUSHT/SHT/U480  ( .ZN(\ALUSHT/pkshtout[14] ), .A(
        \ALUSHT/SHT/n2331 ), .B(\ALUSHT/SHT/n2332 ) );
    snl_oai222x0 \ALUSHT/SHT/U962  ( .ZN(\ALUSHT/SHT/n2762 ), .A(
        \ALUSHT/SHT/n3001 ), .B(\ALUSHT/SHT/n2615 ), .C(\ALUSHT/SHT/n2691 ), 
        .D(\ALUSHT/SHT/n2619 ), .E(\phshtd[1] ), .F(\ALUSHT/SHT/n2692 ) );
    snl_oa2222x1 \ALUSHT/SHT/U1059  ( .Z(\ALUSHT/SHT/n3104 ), .A(
        \ALUSHT/SHT/n3105 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2977 ), 
        .D(\ALUSHT/SHT/n2627 ), .E(\ALUSHT/SHT/n2448 ), .F(\ALUSHT/SHT/n2501 ), 
        .G(\ALUSHT/SHT/n3068 ), .H(\ALUSHT/SHT/n2638 ) );
    snl_invx05 \ALUSHT/SHT/U530  ( .ZN(\ALUSHT/SHT/n2372 ), .A(\poshtfnc[1] )
         );
    snl_invx05 \ALUSHT/SHT/U537  ( .ZN(\ALUSHT/SHT/n2511 ), .A(\pgaluina[13] )
         );
    snl_nand02x1 \ALUSHT/SHT/U600  ( .ZN(\ALUSHT/SHT/n2625 ), .A(
        \ALUSHT/SHT/n2477 ), .B(\ALUSHT/SHT/n2382 ) );
    snl_nand02x1 \ALUSHT/SHT/U607  ( .ZN(\ALUSHT/SHT/n2630 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_oai122x0 \ALUSHT/SHT/U797  ( .ZN(\ALUSHT/SHT/n2825 ), .A(
        \ALUSHT/SHT/n2654 ), .B(\ALUSHT/SHT/n2619 ), .C(\ALUSHT/SHT/n2943 ), 
        .D(\ALUSHT/SHT/n2499 ), .E(\ALUSHT/SHT/n2616 ) );
    snl_oai122x0 \ALUSHT/SHT/U945  ( .ZN(\ALUSHT/SHT/n2755 ), .A(
        \ALUSHT/SHT/n3049 ), .B(\ALUSHT/SHT/n2642 ), .C(\ALUSHT/SHT/n3050 ), 
        .D(\ALUSHT/SHT/n2536 ), .E(\ALUSHT/SHT/n2748 ) );
    snl_nand12x1 \ALUSHT/SHT/U859  ( .ZN(\ALUSHT/SHT/n2622 ), .A(
        \ALUSHT/SHT/n2444 ), .B(\ALUSHT/SHT/n2376 ) );
    snl_aoi022x1 \ALUSHT/SHT/U790  ( .ZN(\ALUSHT/SHT/n2938 ), .A(
        \pgaluina[25] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[24] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_oai122x0 \ALUSHT/SHT/U942  ( .ZN(\ALUSHT/SHT/n2750 ), .A(
        \ALUSHT/SHT/n3005 ), .B(\ALUSHT/SHT/n2614 ), .C(\ALUSHT/SHT/n3006 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n2384 ) );
    snl_nand02x1 \ALUSHT/SHT/U487  ( .ZN(\ALUSHT/pkshtout[21] ), .A(
        \ALUSHT/SHT/n2345 ), .B(\ALUSHT/SHT/n2346 ) );
    snl_oai122x0 \ALUSHT/SHT/U965  ( .ZN(\ALUSHT/SHT/n3058 ), .A(
        \ALUSHT/SHT/n2959 ), .B(\ALUSHT/SHT/n2627 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n3057 ), .E(\ALUSHT/SHT/n2768 ) );
    snl_oai223x0 \ALUSHT/SHT/U517  ( .ZN(\ALUSHT/SHT/n2461 ), .A(\phshtd[0] ), 
        .B(\phshtd[5] ), .C(\ALUSHT/SHT/n2462 ), .D(\ALUSHT/SHT/n2463 ), .E(
        \ALUSHT/SHT/n2464 ), .F(\ALUSHT/SHT/n2465 ), .G(\ALUSHT/SHT/n2466 ) );
    snl_aoi222x0 \ALUSHT/SHT/U328  ( .ZN(\ALUSHT/SHT/n2897 ), .A(
        \ALUSHT/SHT/n2849 ), .B(\ALUSHT/SHT/n2757 ), .C(\ALUSHT/SHT/n2810 ), 
        .D(\ALUSHT/SHT/n2811 ), .E(\ALUSHT/SHT/n2662 ), .F(\ALUSHT/SHT/n2759 )
         );
    snl_aoi2222x0 \ALUSHT/SHT/U354  ( .ZN(\ALUSHT/SHT/n2316 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2738 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2739 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[14] ), 
        .G(\ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2740 ) );
    snl_nand02x2 \ALUSHT/SHT/U368  ( .ZN(\ALUSHT/SHT/n2392 ), .A(
        \ALUSHT/SHT/n2386 ), .B(\ALUSHT/SHT/n2427 ) );
    snl_oai122x0 \ALUSHT/SHT/U579  ( .ZN(\ALUSHT/SHT/n2599 ), .A(
        \ALUSHT/SHT/n2555 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2554 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_nor02x1 \ALUSHT/SHT/U627  ( .ZN(\ALUSHT/SHT/n2444 ), .A(
        \ALUSHT/SHT/n2372 ), .B(\poshtfnc[0] ) );
    snl_oai2222x0 \ALUSHT/SHT/U1079  ( .ZN(\ALUSHT/SHT/n2893 ), .A(
        \ALUSHT/SHT/n3049 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n3051 ), 
        .D(\ALUSHT/SHT/n2627 ), .E(\ALUSHT/SHT/n3050 ), .F(\ALUSHT/SHT/n2638 ), 
        .G(\phshtd[4] ), .H(\ALUSHT/SHT/n2527 ) );
    snl_invx1 \ALUSHT/SHT/U445  ( .ZN(\ALUSHT/SHT/n2492 ), .A(
        \ALUSHT/SHT/n2415 ) );
    snl_invx1 \ALUSHT/SHT/U462  ( .ZN(\ALUSHT/SHT/n2427 ), .A(\phshtd[3] ) );
    snl_nand14x0 \ALUSHT/SHT/U649  ( .ZN(\ALUSHT/SHT/n2703 ), .A(
        \ALUSHT/SHT/n2553 ), .B(\ALUSHT/SHT/n2550 ), .C(\ALUSHT/SHT/n2546 ), 
        .D(\ALUSHT/SHT/n2543 ) );
    snl_oai222x0 \ALUSHT/SHT/U1017  ( .ZN(\ALUSHT/SHT/n2796 ), .A(
        \ALUSHT/SHT/n3018 ), .B(\ALUSHT/SHT/n2615 ), .C(\ALUSHT/SHT/n2689 ), 
        .D(\ALUSHT/SHT/n2619 ), .E(\phshtd[1] ), .F(\ALUSHT/SHT/n3084 ) );
    snl_invx05 \ALUSHT/SHT/U810  ( .ZN(\ALUSHT/SHT/n2951 ), .A(
        \ALUSHT/SHT/n2681 ) );
    snl_aoi122x0 \ALUSHT/SHT/U980  ( .ZN(\ALUSHT/SHT/n3067 ), .A(
        \pgaluina[18] ), .B(\ALUSHT/SHT/n2418 ), .C(\ALUSHT/SHT/n2382 ), .D(
        \ALUSHT/SHT/n2979 ), .E(\ALUSHT/SHT/n2419 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U1030  ( .ZN(\ALUSHT/SHT/n3093 ), .A(
        \ALUSHT/SHT/n2793 ), .B(\ALUSHT/SHT/n2298 ), .C(\ALUSHT/SHT/n2533 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U752  ( .ZN(\ALUSHT/SHT/n2400 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[19] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[20] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[21] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[18] ) );
    snl_invx05 \ALUSHT/SHT/U775  ( .ZN(\ALUSHT/SHT/n2555 ), .A(
        \ALUSHT/SHT/n2863 ) );
    snl_oai2222x0 \ALUSHT/SHT/U837  ( .ZN(\ALUSHT/SHT/n2726 ), .A(
        \ALUSHT/SHT/n2980 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2963 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n2969 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2976 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_nand02x1 \ALUSHT/SHT/U479  ( .ZN(\ALUSHT/pkshtout[13] ), .A(
        \ALUSHT/SHT/n2329 ), .B(\ALUSHT/SHT/n2330 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U749  ( .ZN(\ALUSHT/SHT/n2398 ), .A(
        \ALUSHT/SHT/n2631 ), .B(\pgaluina[27] ), .C(\ALUSHT/SHT/n2541 ), .D(
        \pgaluina[28] ), .E(\ALUSHT/SHT/n2506 ), .F(\pgaluina[29] ), .G(
        \ALUSHT/SHT/n2505 ), .H(\pgaluina[26] ) );
    snl_invx05 \ALUSHT/SHT/U937  ( .ZN(\ALUSHT/SHT/n3049 ), .A(
        \ALUSHT/SHT/n2804 ) );
    snl_oai122x0 \ALUSHT/SHT/U1087  ( .ZN(\ALUSHT/SHT/n2907 ), .A(
        \ALUSHT/SHT/n3016 ), .B(\ALUSHT/SHT/n2454 ), .C(\ALUSHT/SHT/n3002 ), 
        .D(\ALUSHT/SHT/n2642 ), .E(\ALUSHT/SHT/n2905 ) );
    snl_invx05 \ALUSHT/SHT/U1117  ( .ZN(\ALUSHT/SHT/n2597 ), .A(
        \ALUSHT/SHT/n2594 ) );
    snl_bufx1 \ALUSHT/SHT/U373  ( .Z(\ALUSHT/SHT/n2300 ), .A(
        \ALUSHT/SHT/n2615 ) );
    snl_invx05 \ALUSHT/SHT/U545  ( .ZN(\ALUSHT/SHT/n2519 ), .A(\pgaluina[5] )
         );
    snl_oa222x1 \ALUSHT/SHT/U562  ( .Z(\ALUSHT/SHT/n2550 ), .A(
        \ALUSHT/SHT/n2396 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2551 ), 
        .D(\ALUSHT/SHT/n2538 ), .E(\ALUSHT/SHT/n2552 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_nand14x0 \ALUSHT/SHT/U652  ( .ZN(\ALUSHT/SHT/n2706 ), .A(
        \ALUSHT/SHT/n2591 ), .B(\ALUSHT/SHT/n2589 ), .C(\ALUSHT/SHT/n2586 ), 
        .D(\ALUSHT/SHT/n2583 ) );
    snl_aoi012x1 \ALUSHT/SHT/U675  ( .ZN(\ALUSHT/SHT/n2771 ), .A(
        \ALUSHT/SHT/n2423 ), .B(\pgaluina[25] ), .C(\ALUSHT/SHT/n2419 ) );
    snl_oai2222x0 \ALUSHT/SHT/U880  ( .ZN(\ALUSHT/SHT/n2731 ), .A(
        \ALUSHT/SHT/n3009 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2496 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n3016 ), .F(\ALUSHT/SHT/n2642 ), 
        .G(\ALUSHT/SHT/n3014 ), .H(\ALUSHT/SHT/n2454 ) );
    snl_invx05 \ALUSHT/SHT/U910  ( .ZN(\ALUSHT/SHT/n3032 ), .A(
        \ALUSHT/SHT/n2881 ) );
    snl_aoi122x0 \ALUSHT/SHT/U384  ( .ZN(\ALUSHT/SHT/n2333 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[23] ), .C(\ALUSHT/SHT/n2645 ), .D(
        \pgaluina[15] ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U396  ( .ZN(\ALUSHT/SHT/n2332 ), .A(
        \ALUSHT/SHT/n2660 ), .B(\ALUSHT/SHT/n2882 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2883 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[6] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2884 ) );
    snl_aoi2222x2 \ALUSHT/SHT/U417  ( .ZN(\ALUSHT/SHT/n2330 ), .A(
        \ALUSHT/SHT/n2660 ), .B(\ALUSHT/SHT/n2888 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2889 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[5] ), .G(
        \ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2890 ) );
    snl_invx05 \ALUSHT/SHT/U727  ( .ZN(\ALUSHT/SHT/n2438 ), .A(
        \ALUSHT/SHT/n2463 ) );
    snl_oai122x0 \ALUSHT/SHT/U959  ( .ZN(\ALUSHT/SHT/n2757 ), .A(
        \ALUSHT/SHT/n2943 ), .B(\ALUSHT/SHT/n2619 ), .C(\ALUSHT/SHT/n2941 ), 
        .D(\ALUSHT/SHT/n2499 ), .E(\ALUSHT/SHT/n2653 ) );
    snl_aoi2222x0 \ALUSHT/SHT/U1045  ( .ZN(\ALUSHT/SHT/n3099 ), .A(
        \ALUSHT/SHT/n2967 ), .B(\ALUSHT/SHT/n2468 ), .C(\ALUSHT/SHT/n2965 ), 
        .D(\ALUSHT/SHT/n2428 ), .E(\ALUSHT/SHT/n2970 ), .F(\ALUSHT/SHT/n2663 ), 
        .G(\ALUSHT/SHT/n2429 ), .H(\ALUSHT/SHT/n2911 ) );
    snl_oa2222x1 \ALUSHT/SHT/U1062  ( .Z(\ALUSHT/SHT/n3106 ), .A(
        \ALUSHT/SHT/n3107 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2998 ), 
        .D(\ALUSHT/SHT/n2627 ), .E(\ALUSHT/SHT/n3000 ), .F(\ALUSHT/SHT/n2501 ), 
        .G(\ALUSHT/SHT/n3062 ), .H(\ALUSHT/SHT/n2638 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U865  ( .ZN(\ALUSHT/SHT/n3005 ), .A(
        \pgaluina[31] ), .B(\ALUSHT/SHT/n2910 ), .C(\ALUSHT/SHT/n2917 ) );
    snl_nand02x3 \ALUSHT/SHT/U405  ( .ZN(\ALUSHT/SHT/n2502 ), .A(\phshtd[4] ), 
        .B(\ALUSHT/SHT/n2441 ) );
    snl_aoi012x4 \ALUSHT/SHT/U430  ( .ZN(\ALUSHT/SHT/n2693 ), .A(
        \ALUSHT/SHT/n2694 ), .B(\ALUSHT/SHT/n2695 ), .C(\ALUSHT/SHT/n2696 ) );
    snl_oai122x0 \ALUSHT/SHT/U587  ( .ZN(\ALUSHT/SHT/n2607 ), .A(
        \ALUSHT/SHT/n2582 ), .B(\ALUSHT/SHT/n2510 ), .C(\ALUSHT/SHT/n2387 ), 
        .D(\ALUSHT/SHT/n2502 ), .E(\ALUSHT/SHT/n2594 ) );
    snl_aoi012x1 \ALUSHT/SHT/U842  ( .ZN(\ALUSHT/SHT/n2987 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[29] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_nand02x1 \ALUSHT/SHT/U595  ( .ZN(\ALUSHT/SHT/n2451 ), .A(
        \ALUSHT/SHT/n2298 ), .B(\ALUSHT/SHT/n2498 ) );
    snl_aoi222x0 \ALUSHT/SHT/U690  ( .ZN(\ALUSHT/SHT/n2346 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2844 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2845 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2841 )
         );
    snl_aoi122x0 \ALUSHT/SHT/U700  ( .ZN(\ALUSHT/SHT/n2304 ), .A(
        \ALUSHT/SHT/n2634 ), .B(\pgaluina[8] ), .C(\ALUSHT/SHT/n2643 ), .D(
        \ALUSHT/SHT/n2907 ), .E(\ALUSHT/SHT/n2906 ) );
    snl_invx05 \ALUSHT/SHT/U735  ( .ZN(\ALUSHT/SHT/n2565 ), .A(
        \ALUSHT/SHT/n2394 ) );
    snl_aoi122x2 \ALUSHT/SHT/U422  ( .ZN(\ALUSHT/SHT/n2359 ), .A(
        \ALUSHT/SHT/n2644 ), .B(\pgaluina[4] ), .C(\pgaluina[28] ), .D(
        \ALUSHT/SHT/n2788 ), .E(\ALUSHT/SHT/n2367 ) );
    snl_aoi022x1 \ALUSHT/SHT/U877  ( .ZN(\ALUSHT/SHT/n3015 ), .A(
        \pgaluina[16] ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[15] ), .D(
        \ALUSHT/SHT/n2910 ) );
    snl_aoi222x0 \ALUSHT/SHT/U682  ( .ZN(\ALUSHT/SHT/n2362 ), .A(
        \ALUSHT/SHT/n2643 ), .B(\ALUSHT/SHT/n2802 ), .C(\ALUSHT/SHT/n2639 ), 
        .D(\ALUSHT/SHT/n2803 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2787 )
         );
    snl_nor02x1 \ALUSHT/SHT/U712  ( .ZN(\ALUSHT/SHT/n2410 ), .A(
        \ALUSHT/SHT/n2626 ), .B(\ALUSHT/SHT/n2382 ) );
    snl_aoi012x1 \ALUSHT/SHT/U850  ( .ZN(\ALUSHT/SHT/n2412 ), .A(
        \ALUSHT/SHT/n2491 ), .B(\pgaluina[19] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1057  ( .ZN(\ALUSHT/SHT/n2859 ), .A(
        \ALUSHT/SHT/n3103 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3096 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3098 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3100 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_oai2222x0 \ALUSHT/SHT/U1070  ( .ZN(\ALUSHT/SHT/n2884 ), .A(
        \ALUSHT/SHT/n2969 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n3102 ), 
        .D(\ALUSHT/SHT/n2300 ), .E(\ALUSHT/SHT/n3104 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n2963 ), .H(\ALUSHT/SHT/n2299 ) );
    snl_aoi222x0 \ALUSHT/SHT/U333  ( .ZN(\ALUSHT/SHT/n2692 ), .A(
        \ALUSHT/SHT/n2994 ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2411 ), 
        .D(\ALUSHT/SHT/n2539 ), .E(\ALUSHT/SHT/n3027 ), .F(\phshtd[2] ) );
    snl_aoi2222x0 \ALUSHT/SHT/U346  ( .ZN(\ALUSHT/SHT/n2334 ), .A(
        \ALUSHT/SHT/n2634 ), .B(\pgaluina[7] ), .C(\ALUSHT/SHT/n2639 ), .D(
        \ALUSHT/SHT/n2878 ), .E(\ALUSHT/SHT/n2641 ), .F(\ALUSHT/SHT/n2875 ), 
        .G(\ALUSHT/SHT/n2643 ), .H(\ALUSHT/SHT/n2879 ) );
    snl_invx05 \ALUSHT/SHT/U539  ( .ZN(\ALUSHT/SHT/n2513 ), .A(\pgaluina[11] )
         );
    snl_oa022x1 \ALUSHT/SHT/U557  ( .Z(\ALUSHT/SHT/n2535 ), .A(
        \ALUSHT/SHT/n2529 ), .B(\ALUSHT/SHT/n2392 ), .C(\ALUSHT/SHT/n2385 ), 
        .D(\ALUSHT/SHT/n2399 ) );
    snl_nor03x0 \ALUSHT/SHT/U609  ( .ZN(\ALUSHT/SHT/n2633 ), .A(\poshtfnc[1] ), 
        .B(\poshtfnc[2] ), .C(\ALUSHT/SHT/n2623 ) );
    snl_oai2222x0 \ALUSHT/SHT/U799  ( .ZN(\ALUSHT/SHT/n2727 ), .A(
        \ALUSHT/SHT/n2937 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2493 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2944 ), .F(\ALUSHT/SHT/n2642 ), 
        .G(\ALUSHT/SHT/n2942 ), .H(\ALUSHT/SHT/n2454 ) );
    snl_oa222x1 \ALUSHT/SHT/U1039  ( .Z(\ALUSHT/SHT/n3097 ), .A(
        \ALUSHT/SHT/n2959 ), .B(\ALUSHT/SHT/n2640 ), .C(\ALUSHT/SHT/n2961 ), 
        .D(\ALUSHT/SHT/n2501 ), .E(\ALUSHT/SHT/n3057 ), .F(\ALUSHT/SHT/n2427 )
         );
    snl_aoi2222x0 \ALUSHT/SHT/U361  ( .ZN(\ALUSHT/SHT/n2308 ), .A(
        \ALUSHT/SHT/n2721 ), .B(\ALUSHT/SHT/n2794 ), .C(\ALUSHT/SHT/n2723 ), 
        .D(\ALUSHT/SHT/n2795 ), .E(\ALUSHT/SHT/n2634 ), .F(\pgaluina[10] ), 
        .G(\ALUSHT/SHT/n2639 ), .H(\ALUSHT/SHT/n2796 ) );
    snl_muxi21x1 \ALUSHT/SHT/U640  ( .ZN(\ALUSHT/SHT/n2375 ), .A(
        \ALUSHT/SHT/n2665 ), .B(\ALUSHT/SHT/n2666 ), .S(\ALUSHT/SHT/n2383 ) );
    snl_aoi012x1 \ALUSHT/SHT/U667  ( .ZN(\ALUSHT/SHT/n2732 ), .A(
        \ALUSHT/SHT/n2651 ), .B(\pgaluina[7] ), .C(\ALUSHT/SHT/n2492 ) );
    snl_oai222x0 \ALUSHT/SHT/U925  ( .ZN(\ALUSHT/SHT/n2743 ), .A(
        \ALUSHT/SHT/n3041 ), .B(\ALUSHT/SHT/n2451 ), .C(\ALUSHT/SHT/n2406 ), 
        .D(\ALUSHT/SHT/n2380 ), .E(\ALUSHT/SHT/n3042 ), .F(\ALUSHT/SHT/n2454 )
         );
    snl_aoi222x1 \ALUSHT/SHT/U457  ( .ZN(\ALUSHT/SHT/n2828 ), .A(
        \ALUSHT/SHT/n2548 ), .B(\ALUSHT/SHT/n2829 ), .C(\ALUSHT/SHT/n2659 ), 
        .D(\ALUSHT/SHT/n2830 ), .E(\ALUSHT/SHT/n2810 ), .F(\ALUSHT/SHT/n2831 )
         );
    snl_nand02x1 \ALUSHT/SHT/U470  ( .ZN(\ALUSHT/pkshtout[4] ), .A(
        \ALUSHT/SHT/n2311 ), .B(\ALUSHT/SHT/n2312 ) );
    snl_oa222x1 \ALUSHT/SHT/U570  ( .Z(\ALUSHT/SHT/n2578 ), .A(
        \ALUSHT/SHT/n2579 ), .B(\ALUSHT/SHT/n2380 ), .C(\ALUSHT/SHT/n2534 ), 
        .D(\ALUSHT/SHT/n2510 ), .E(\ALUSHT/SHT/n2580 ), .F(\ALUSHT/SHT/n2502 )
         );
    snl_nand02x1 \ALUSHT/SHT/U819  ( .ZN(\ALUSHT/SHT/n2491 ), .A(\phshtd[5] ), 
        .B(\ALUSHT/SHT/n2374 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U892  ( .ZN(\ALUSHT/SHT/n3022 ), .A(
        \ALUSHT/SHT/n2877 ), .B(\ALUSHT/SHT/n2298 ), .C(\ALUSHT/SHT/n2573 ) );
    snl_invx05 \ALUSHT/SHT/U902  ( .ZN(\ALUSHT/SHT/n3029 ), .A(
        \ALUSHT/SHT/n2783 ) );
    snl_invx05 \ALUSHT/SHT/U1122  ( .ZN(\ALUSHT/SHT/n2453 ), .A(
        \ALUSHT/SHT/n2495 ) );
    snl_oai113x0 \ALUSHT/SHT/U989  ( .ZN(\ALUSHT/SHT/n2439 ), .A(
        \ALUSHT/SHT/n2625 ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2512 ), 
        .D(\ALUSHT/SHT/n2916 ), .E(\ALUSHT/SHT/n2777 ) );
    snl_aoi022x1 \ALUSHT/SHT/U1095  ( .ZN(\ALUSHT/SHT/n2440 ), .A(
        \ALUSHT/SHT/n3075 ), .B(\ALUSHT/SHT/n2504 ), .C(\ALUSHT/SHT/n2680 ), 
        .D(\phshtd[0] ) );
    snl_invx05 \ALUSHT/SHT/U1105  ( .ZN(\ALUSHT/SHT/n3089 ), .A(
        \ALUSHT/SHT/n2972 ) );
    snl_invx05 \ALUSHT/SHT/U740  ( .ZN(\ALUSHT/SHT/n2791 ), .A(
        \ALUSHT/SHT/n2538 ) );
    snl_oai012x1 \ALUSHT/SHT/U802  ( .ZN(\ALUSHT/SHT/n2778 ), .A(
        \ALUSHT/SHT/n2520 ), .B(\ALUSHT/SHT/n2625 ), .C(\ALUSHT/SHT/n2916 ) );
    snl_oai113x0 \ALUSHT/SHT/U992  ( .ZN(\ALUSHT/SHT/n3073 ), .A(
        \ALUSHT/SHT/n2625 ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2513 ), 
        .D(\ALUSHT/SHT/n2916 ), .E(\ALUSHT/SHT/n2774 ) );
    snl_oa122x1 \ALUSHT/SHT/U767  ( .Z(\ALUSHT/SHT/n2561 ), .A(
        \ALUSHT/SHT/n2923 ), .B(\ALUSHT/SHT/n2388 ), .C(\ALUSHT/SHT/n2587 ), 
        .D(\ALUSHT/SHT/n2399 ), .E(\ALUSHT/SHT/n2699 ) );
    snl_nand02x1 \ALUSHT/SHT/U612  ( .ZN(\ALUSHT/SHT/n2636 ), .A(
        \ALUSHT/SHT/n2477 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U782  ( .ZN(\ALUSHT/SHT/n2456 ), .A(
        \ALUSHT/SHT/n2386 ), .B(\ALUSHT/SHT/n2407 ), .C(\ALUSHT/SHT/n2616 ) );
    snl_oai012x1 \ALUSHT/SHT/U825  ( .ZN(\ALUSHT/SHT/n2965 ), .A(
        \ALUSHT/SHT/n2652 ), .B(\ALUSHT/SHT/n2397 ), .C(\ALUSHT/SHT/n2415 ) );
    snl_oai222x0 \ALUSHT/SHT/U889  ( .ZN(\ALUSHT/SHT/n2733 ), .A(
        \ALUSHT/SHT/n3020 ), .B(\ALUSHT/SHT/n2454 ), .C(\ALUSHT/SHT/n3019 ), 
        .D(\ALUSHT/SHT/n2451 ), .E(\ALUSHT/SHT/n2573 ), .F(\ALUSHT/SHT/n2380 )
         );
    snl_invx05 \ALUSHT/SHT/U919  ( .ZN(\ALUSHT/SHT/n3040 ), .A(
        \ALUSHT/SHT/n3039 ) );
    snl_invx05 \ALUSHT/SHT/U1005  ( .ZN(\ALUSHT/SHT/n3079 ), .A(
        \ALUSHT/SHT/n2861 ) );
    snl_aoi0b12x0 \ALUSHT/SHT/U1022  ( .ZN(\ALUSHT/SHT/n3087 ), .A(
        \ALUSHT/SHT/n2750 ), .B(\ALUSHT/SHT/n2298 ), .C(\ALUSHT/SHT/n2527 ) );
    snl_nor02x1 \ALUSHT/SHT/U505  ( .ZN(\ALUSHT/SHT/n2394 ), .A(
        \ALUSHT/SHT/n2392 ), .B(\ALUSHT/SHT/n2395 ) );
    snl_aoi022x1 \ALUSHT/SHT/U522  ( .ZN(\ALUSHT/SHT/n2487 ), .A(
        \ALUSHT/SHT/n2468 ), .B(\ALUSHT/SHT/n2488 ), .C(\ALUSHT/SHT/n2298 ), 
        .D(\ALUSHT/SHT/n2489 ) );
    snl_oai2222x0 \ALUSHT/SHT/U950  ( .ZN(\ALUSHT/SHT/n2754 ), .A(
        \ALUSHT/SHT/n2689 ), .B(\ALUSHT/SHT/n2302 ), .C(\ALUSHT/SHT/n2980 ), 
        .D(\ALUSHT/SHT/n2615 ), .E(\ALUSHT/SHT/n3018 ), .F(\ALUSHT/SHT/n2301 ), 
        .G(\ALUSHT/SHT/n3040 ), .H(\ALUSHT/SHT/n2619 ) );
    snl_aoi022x1 \ALUSHT/SHT/U314  ( .ZN(\ALUSHT/SHT/n2672 ), .A(\pgaluina[2] 
        ), .B(\ALUSHT/SHT/n2650 ), .C(\pgaluina[1] ), .D(\ALUSHT/SHT/n2910 )
         );
    snl_nand02x1 \ALUSHT/SHT/U495  ( .ZN(\ALUSHT/pkshtout[29] ), .A(
        \ALUSHT/SHT/n2361 ), .B(\ALUSHT/SHT/n2362 ) );
    snl_aoi122x2 \ALUSHT/SHT/U439  ( .ZN(\ALUSHT/SHT/n2572 ), .A(
        \ALUSHT/SHT/n2584 ), .B(\ALUSHT/SHT/n2694 ), .C(\ALUSHT/SHT/n2698 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2914 ) );
    snl_nor02x1 \ALUSHT/SHT/U635  ( .ZN(\ALUSHT/SHT/n2659 ), .A(
        \ALUSHT/SHT/n2382 ), .B(\ALUSHT/SHT/n2441 ) );
    snl_aoi222x0 \ALUSHT/SHT/U977  ( .ZN(\ALUSHT/SHT/n2679 ), .A(
        \ALUSHT/SHT/n3063 ), .B(\ALUSHT/SHT/n2404 ), .C(\ALUSHT/SHT/n2420 ), 
        .D(\ALUSHT/SHT/n2390 ), .E(\ALUSHT/SHT/n2386 ), .F(\ALUSHT/SHT/n3065 )
         );
    snl_oai022x1 \ALUSHT/SHT/U699  ( .ZN(\ALUSHT/SHT/n2906 ), .A(
        \ALUSHT/SHT/n2482 ), .B(\ALUSHT/SHT/n2632 ), .C(\ALUSHT/SHT/n2476 ), 
        .D(\ALUSHT/SHT/n2621 ) );
    snl_invx05 \ALUSHT/SHT/U709  ( .ZN(\ALUSHT/SHT/n2539 ), .A(
        \ALUSHT/SHT/n2392 ) );
    snl_nand12x1 \REG_2/ph8dec_2/U6  ( .ZN(\REG_2/ncnt2[2] ), .A(ph_byrtendh), 
        .B(\REG_2/ph8dec_2/n20 ) );
    snl_invx05 \REG_2/ph8dec_2/U7  ( .ZN(\REG_2/ncnt2[0] ), .A(
        \REG_2/RETCNT[3] ) );
    snl_aoi022x1 \REG_2/ph8dec_2/U8  ( .ZN(\REG_2/ncnt2[1] ), .A(
        \REG_2/RETCNT[4] ), .B(\REG_2/ncnt2[0] ), .C(\REG_2/ph8dec_2/n21 ), 
        .D(\REG_2/RETCNT[3] ) );
    snl_nor03x0 \REG_2/ph8dec_2/U9  ( .ZN(ph_byrtendh), .A(\REG_2/RETCNT[3] ), 
        .B(\REG_2/RETCNT[5] ), .C(\REG_2/RETCNT[4] ) );
    snl_oai012x1 \REG_2/ph8dec_2/U10  ( .ZN(\REG_2/ph8dec_2/n20 ), .A(
        \REG_2/RETCNT[4] ), .B(\REG_2/RETCNT[3] ), .C(\REG_2/RETCNT[5] ) );
    snl_invx05 \REG_2/ph8dec_2/U11  ( .ZN(\REG_2/ph8dec_2/n21 ), .A(
        \REG_2/RETCNT[4] ) );
    snl_invx1 \CODEQ/phque34_1/U8  ( .ZN(\CODEQ/phque34_1/n753 ), .A(
        \CODEQ/phque34_1/n761 ) );
    snl_and02x2 \CODEQ/phque34_1/U13  ( .Z(\CODEQ/phque34_1/n757 ), .A(
        ph_exe_ah), .B(ph_exe_ch) );
    snl_muxi21x2 \CODEQ/phque34_1/U14  ( .ZN(\CODEQ/phque34_1/n759 ), .A(
        \CODEQ/phque34_1/n761 ), .B(\CODEQ/phque34_1/n762 ), .S(
        \CODEQ/phque34_1/n763 ) );
    snl_oai022x1 \CODEQ/phque34_1/U21  ( .ZN(\stream4[5] ), .A(
        \CODEQ/nqueue1[5] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[5] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U54  ( .ZN(\stream4[38] ), .A(
        \CODEQ/nqueue1[38] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[38] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U73  ( .ZN(\stream4[57] ), .A(
        \CODEQ/nqueue1[57] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[57] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U113  ( .ZN(\CODEQ/phque34_1/stream3[37] ), 
        .A(\CODEQ/nqueue2[37] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[37] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U134  ( .ZN(\stream3[58] ), .A(
        \CODEQ/nqueue2[58] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[58] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U96  ( .ZN(\stream3[20] ), .A(
        \CODEQ/nqueue1[20] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[20] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U68  ( .ZN(\stream4[52] ), .A(
        \CODEQ/nqueue1[52] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[52] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U108  ( .ZN(\stream3[32] ), .A(
        \CODEQ/nqueue1[32] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[32] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_nand02x1 \CODEQ/phque34_1/U141  ( .ZN(\CODEQ/phque34_1/n765 ), .A(
        ph_exe_bh), .B(ph_exe_dh) );
    snl_oai022x1 \CODEQ/phque34_1/U28  ( .ZN(\stream4[12] ), .A(
        \CODEQ/nqueue1[12] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[12] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U33  ( .ZN(\stream4[17] ), .A(
        \CODEQ/nqueue1[17] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[17] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U34  ( .ZN(\stream4[18] ), .A(
        \CODEQ/nqueue1[18] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[18] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U41  ( .ZN(\stream4[25] ), .A(
        \CODEQ/nqueue1[25] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[25] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U46  ( .ZN(\stream4[30] ), .A(
        \CODEQ/nqueue1[30] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[30] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U61  ( .ZN(\stream4[45] ), .A(
        \CODEQ/nqueue1[45] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[45] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U84  ( .ZN(\stream3[8] ), .A(
        \CODEQ/nqueue2[8] ), .B(\CODEQ/phque34_1/n755 ), .C(\CODEQ/nqueue1[8] 
        ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U101  ( .ZN(\stream3[25] ), .A(
        \CODEQ/nqueue2[25] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[25] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U126  ( .ZN(\stream3[50] ), .A(
        \CODEQ/nqueue2[50] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[50] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U66  ( .ZN(\stream4[50] ), .A(
        \CODEQ/nqueue1[50] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[50] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U106  ( .ZN(\stream3[30] ), .A(
        \CODEQ/nqueue2[30] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[30] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U121  ( .ZN(\stream3[45] ), .A(
        \CODEQ/nqueue2[45] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[45] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U83  ( .ZN(\stream3[7] ), .A(
        \CODEQ/nqueue2[7] ), .B(\CODEQ/phque34_1/n760 ), .C(\CODEQ/nqueue1[7] 
        ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U98  ( .ZN(\stream3[22] ), .A(
        \CODEQ/nqueue1[22] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[22] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U26  ( .ZN(\stream4[10] ), .A(
        \CODEQ/nqueue1[10] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[10] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U48  ( .ZN(\stream4[32] ), .A(
        \CODEQ/nqueue1[32] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[32] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U128  ( .ZN(\stream3[52] ), .A(
        \CODEQ/nqueue1[52] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[52] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_bufx1 \CODEQ/phque34_1/U9  ( .Z(\CODEQ/phque34_1/n754 ), .A(
        \CODEQ/phque34_1/n758 ) );
    snl_bufx1 \CODEQ/phque34_1/U12  ( .Z(\CODEQ/phque34_1/n756 ), .A(
        \CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U35  ( .ZN(\stream4[19] ), .A(
        \CODEQ/nqueue1[19] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[19] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U53  ( .ZN(\stream4[37] ), .A(
        \CODEQ/nqueue1[37] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[37] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U91  ( .ZN(\stream3[15] ), .A(
        \CODEQ/nqueue1[15] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[15] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U74  ( .ZN(\stream4[58] ), .A(
        \CODEQ/nqueue1[58] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[58] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U114  ( .ZN(\CODEQ/phque34_1/stream3[38] ), 
        .A(\CODEQ/nqueue2[38] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[38] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U133  ( .ZN(\stream3[57] ), .A(
        \CODEQ/nqueue2[57] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[57] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U99  ( .ZN(\stream3[23] ), .A(
        \CODEQ/nqueue2[23] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[23] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U27  ( .ZN(\stream4[11] ), .A(
        \CODEQ/nqueue1[11] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[11] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U40  ( .ZN(\stream4[24] ), .A(
        \CODEQ/nqueue1[24] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[24] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U82  ( .ZN(\stream3[6] ), .A(
        \CODEQ/nqueue1[6] ), .B(\CODEQ/phque34_1/n759 ), .C(\CODEQ/nqueue2[6] 
        ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U52  ( .ZN(\stream4[36] ), .A(
        \CODEQ/nqueue1[36] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[36] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U67  ( .ZN(\stream4[51] ), .A(
        \CODEQ/nqueue1[51] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[51] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U107  ( .ZN(\stream3[31] ), .A(
        \CODEQ/nqueue1[31] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[31] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U120  ( .ZN(\stream3[44] ), .A(
        \CODEQ/nqueue1[44] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[44] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U75  ( .ZN(\stream4[59] ), .A(
        \CODEQ/nqueue1[59] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[59] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U115  ( .ZN(\CODEQ/phque34_1/stream3[39] ), 
        .A(\CODEQ/nqueue2[39] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[39] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U132  ( .ZN(\stream3[56] ), .A(
        \CODEQ/nqueue1[56] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[56] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U90  ( .ZN(\stream3[14] ), .A(
        \CODEQ/nqueue1[14] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[14] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_bufx1 \CODEQ/phque34_1/U10  ( .Z(\CODEQ/phque34_1/n755 ), .A(
        \CODEQ/phque34_1/n760 ) );
    snl_aob1b12x2 \CODEQ/phque34_1/U15  ( .Z(\CODEQ/phque34_1/n758 ), .A(
        ph_exe_dh), .B(ph_exe_bh), .C(ph_exe_ch), .D(ph_exe_ah) );
    snl_oai022x1 \CODEQ/phque34_1/U20  ( .ZN(\stream4[4] ), .A(
        \CODEQ/nqueue1[4] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[4] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U49  ( .ZN(\stream4[33] ), .A(
        \CODEQ/nqueue1[33] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[33] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U129  ( .ZN(\stream3[53] ), .A(
        \CODEQ/nqueue2[53] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[53] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U69  ( .ZN(\stream4[53] ), .A(
        \CODEQ/nqueue1[53] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[53] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U109  ( .ZN(\stream3[33] ), .A(
        \CODEQ/nqueue1[33] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[33] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U29  ( .ZN(\stream4[13] ), .A(
        \CODEQ/nqueue1[13] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[13] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U47  ( .ZN(\stream4[31] ), .A(
        \CODEQ/nqueue1[31] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[31] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U55  ( .ZN(\stream4[39] ), .A(
        \CODEQ/nqueue1[39] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[39] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U72  ( .ZN(\stream4[56] ), .A(
        \CODEQ/nqueue1[56] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[56] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U97  ( .ZN(\stream3[21] ), .A(
        \CODEQ/nqueue1[21] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[21] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_nand02x1 \CODEQ/phque34_1/U140  ( .ZN(\CODEQ/phque34_1/n766 ), .A(
        ph_dec_dh), .B(ph_dec_bh) );
    snl_oai022x1 \CODEQ/phque34_1/U112  ( .ZN(\CODEQ/phque34_1/stream3[36] ), 
        .A(\CODEQ/nqueue1[36] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[36] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U135  ( .ZN(\stream3[59] ), .A(
        \CODEQ/nqueue1[59] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[59] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U60  ( .ZN(\stream4[44] ), .A(
        \CODEQ/nqueue1[44] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[44] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U100  ( .ZN(\stream3[24] ), .A(
        \CODEQ/nqueue1[24] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[24] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U127  ( .ZN(\stream3[51] ), .A(
        \CODEQ/nqueue2[51] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[51] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U85  ( .ZN(\stream3[9] ), .A(
        \CODEQ/nqueue1[9] ), .B(\CODEQ/phque34_1/n759 ), .C(\CODEQ/nqueue2[9] 
        ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U17  ( .ZN(\stream4[1] ), .A(
        \CODEQ/nqueue1[1] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[1] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U22  ( .ZN(\stream4[6] ), .A(
        \CODEQ/nqueue1[6] ), .B(\CODEQ/phque34_1/n753 ), .C(\CODEQ/nqueue2[6] 
        ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U32  ( .ZN(\stream4[16] ), .A(
        \CODEQ/nqueue1[16] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[16] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U39  ( .ZN(\stream4[23] ), .A(
        \CODEQ/nqueue1[23] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[23] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U57  ( .ZN(\stream4[41] ), .A(
        \CODEQ/nqueue1[41] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[41] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_nand02x1 \CODEQ/phque34_1/U137  ( .ZN(\CODEQ/phque34_1/n761 ), .A(
        ph_exe_ah), .B(ph_exe_ch) );
    snl_oai022x1 \CODEQ/phque34_1/U70  ( .ZN(\stream4[54] ), .A(
        \CODEQ/nqueue1[54] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[54] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U110  ( .ZN(\stream3[34] ), .A(
        \CODEQ/nqueue2[34] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[34] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U95  ( .ZN(\stream3[19] ), .A(
        \CODEQ/nqueue1[19] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[19] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U30  ( .ZN(\stream4[14] ), .A(
        \CODEQ/nqueue1[14] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[14] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U79  ( .ZN(\stream3[3] ), .A(
        \CODEQ/nqueue2[3] ), .B(\CODEQ/phque34_1/n760 ), .C(\CODEQ/nqueue1[3] 
        ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U119  ( .ZN(\stream3[43] ), .A(
        \CODEQ/nqueue2[43] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[43] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U42  ( .ZN(\stream4[26] ), .A(
        \CODEQ/nqueue1[26] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[26] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U45  ( .ZN(\stream4[29] ), .A(
        \CODEQ/nqueue1[29] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[29] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U87  ( .ZN(\stream3[11] ), .A(
        \CODEQ/nqueue2[11] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[11] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U125  ( .ZN(\stream3[49] ), .A(
        \CODEQ/nqueue2[49] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[49] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U62  ( .ZN(\stream4[46] ), .A(
        \CODEQ/nqueue1[46] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[46] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U65  ( .ZN(\stream4[49] ), .A(
        \CODEQ/nqueue1[49] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[49] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U102  ( .ZN(\stream3[26] ), .A(
        \CODEQ/nqueue2[26] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[26] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U105  ( .ZN(\stream3[29] ), .A(
        \CODEQ/nqueue2[29] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[29] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U80  ( .ZN(\stream3[4] ), .A(
        \CODEQ/nqueue1[4] ), .B(\CODEQ/phque34_1/n759 ), .C(\CODEQ/nqueue2[4] 
        ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U122  ( .ZN(\stream3[46] ), .A(
        \CODEQ/nqueue1[46] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[46] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_nand12x2 \CODEQ/phque34_1/U11  ( .ZN(\CODEQ/phque34_1/n760 ), .A(
        \CODEQ/phque34_1/n764 ), .B(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U19  ( .ZN(\stream4[3] ), .A(
        \CODEQ/nqueue1[3] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[3] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U25  ( .ZN(\stream4[9] ), .A(
        \CODEQ/nqueue1[9] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[9] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U37  ( .ZN(\stream4[21] ), .A(
        \CODEQ/nqueue1[21] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[21] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U59  ( .ZN(\stream4[43] ), .A(
        \CODEQ/nqueue1[43] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[43] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_nor03x0 \CODEQ/phque34_1/U139  ( .ZN(\CODEQ/phque34_1/n763 ), .A(
        ph_exstgb_h), .B(ph_exstga_h), .C(stage_b) );
    snl_oai022x1 \CODEQ/phque34_1/U89  ( .ZN(\stream3[13] ), .A(
        \CODEQ/nqueue1[13] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[13] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U50  ( .ZN(\stream4[34] ), .A(
        \CODEQ/nqueue1[34] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[34] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U77  ( .ZN(\stream3[1] ), .A(
        \CODEQ/nqueue2[1] ), .B(\CODEQ/phque34_1/n760 ), .C(\CODEQ/nqueue1[1] 
        ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U92  ( .ZN(\stream3[16] ), .A(
        \CODEQ/nqueue2[16] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[16] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U117  ( .ZN(\stream3[41] ), .A(
        \CODEQ/nqueue2[41] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[41] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U58  ( .ZN(\stream4[42] ), .A(
        \CODEQ/nqueue1[42] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[42] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U130  ( .ZN(\stream3[54] ), .A(
        \CODEQ/nqueue1[54] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[54] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_muxi21x1 \CODEQ/phque34_1/U138  ( .ZN(\CODEQ/phque34_1/n764 ), .A(
        \CODEQ/phque34_1/n765 ), .B(\CODEQ/phque34_1/n766 ), .S(
        \CODEQ/phque34_1/n763 ) );
    snl_oai022x1 \CODEQ/phque34_1/U16  ( .ZN(\stream4[0] ), .A(
        \CODEQ/nqueue1[0] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[0] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U18  ( .ZN(\stream4[2] ), .A(
        \CODEQ/nqueue1[2] ), .B(\CODEQ/phque34_1/n753 ), .C(\CODEQ/nqueue2[2] 
        ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U36  ( .ZN(\stream4[20] ), .A(
        \CODEQ/nqueue1[20] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[20] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U43  ( .ZN(\stream4[27] ), .A(
        \CODEQ/nqueue1[27] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[27] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U64  ( .ZN(\stream4[48] ), .A(
        \CODEQ/nqueue1[48] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[48] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U81  ( .ZN(\stream3[5] ), .A(
        \CODEQ/nqueue2[5] ), .B(\CODEQ/phque34_1/n760 ), .C(\CODEQ/nqueue1[5] 
        ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U104  ( .ZN(\stream3[28] ), .A(
        \CODEQ/nqueue1[28] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[28] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U51  ( .ZN(\stream4[35] ), .A(
        \CODEQ/nqueue1[35] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[35] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U76  ( .ZN(\stream3[0] ), .A(
        \CODEQ/nqueue1[0] ), .B(\CODEQ/phque34_1/n759 ), .C(\CODEQ/nqueue2[0] 
        ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U116  ( .ZN(\stream3[40] ), .A(
        \CODEQ/nqueue2[40] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[40] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U123  ( .ZN(\stream3[47] ), .A(
        \CODEQ/nqueue1[47] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[47] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U131  ( .ZN(\stream3[55] ), .A(
        \CODEQ/nqueue2[55] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[55] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U23  ( .ZN(\stream4[7] ), .A(
        \CODEQ/nqueue1[7] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[7] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U24  ( .ZN(\stream4[8] ), .A(
        \CODEQ/nqueue1[8] ), .B(\CODEQ/phque34_1/n757 ), .C(\CODEQ/nqueue2[8] 
        ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U88  ( .ZN(\stream3[12] ), .A(
        \CODEQ/nqueue1[12] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[12] ), .D(\CODEQ/phque34_1/n755 ) );
    snl_oai022x1 \CODEQ/phque34_1/U93  ( .ZN(\stream3[17] ), .A(
        \CODEQ/nqueue2[17] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[17] ), .D(\CODEQ/phque34_1/n756 ) );
    snl_oai022x1 \CODEQ/phque34_1/U31  ( .ZN(\stream4[15] ), .A(
        \CODEQ/nqueue1[15] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[15] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U38  ( .ZN(\stream4[22] ), .A(
        \CODEQ/nqueue1[22] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[22] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U44  ( .ZN(\stream4[28] ), .A(
        \CODEQ/nqueue1[28] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[28] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U56  ( .ZN(\stream4[40] ), .A(
        \CODEQ/nqueue1[40] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[40] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U94  ( .ZN(\stream3[18] ), .A(
        \CODEQ/nqueue2[18] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[18] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_nand02x1 \CODEQ/phque34_1/U136  ( .ZN(\CODEQ/phque34_1/n762 ), .A(
        ph_dec_ch), .B(ph_dec_ah) );
    snl_oai022x1 \CODEQ/phque34_1/U71  ( .ZN(\stream4[55] ), .A(
        \CODEQ/nqueue1[55] ), .B(\CODEQ/phque34_1/n753 ), .C(
        \CODEQ/nqueue2[55] ), .D(\CODEQ/phque34_1/n754 ) );
    snl_oai022x1 \CODEQ/phque34_1/U111  ( .ZN(\CODEQ/phque34_1/stream3[35] ), 
        .A(\CODEQ/nqueue2[35] ), .B(\CODEQ/phque34_1/n760 ), .C(
        \CODEQ/nqueue1[35] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U124  ( .ZN(\stream3[48] ), .A(
        \CODEQ/nqueue2[48] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[48] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U63  ( .ZN(\stream4[47] ), .A(
        \CODEQ/nqueue1[47] ), .B(\CODEQ/phque34_1/n757 ), .C(
        \CODEQ/nqueue2[47] ), .D(\CODEQ/phque34_1/n758 ) );
    snl_oai022x1 \CODEQ/phque34_1/U86  ( .ZN(\stream3[10] ), .A(
        \CODEQ/nqueue2[10] ), .B(\CODEQ/phque34_1/n755 ), .C(
        \CODEQ/nqueue1[10] ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U103  ( .ZN(\stream3[27] ), .A(
        \CODEQ/nqueue1[27] ), .B(\CODEQ/phque34_1/n756 ), .C(
        \CODEQ/nqueue2[27] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_oai022x1 \CODEQ/phque34_1/U78  ( .ZN(\stream3[2] ), .A(
        \CODEQ/nqueue2[2] ), .B(\CODEQ/phque34_1/n755 ), .C(\CODEQ/nqueue1[2] 
        ), .D(\CODEQ/phque34_1/n759 ) );
    snl_oai022x1 \CODEQ/phque34_1/U118  ( .ZN(\stream3[42] ), .A(
        \CODEQ/nqueue1[42] ), .B(\CODEQ/phque34_1/n759 ), .C(
        \CODEQ/nqueue2[42] ), .D(\CODEQ/phque34_1/n760 ) );
    snl_and02x1 \LBUS/ldoecnt_3/U8  ( .Z(ph_ldaoutenh3), .A(ph_lbwrh), .B(
        \LBUS/temp[3] ) );
    snl_nand14x0 \MCD/rd_wt_1/U88  ( .ZN(saenabl1), .A(rrmw1), .B(
        \MCD/rd_wt_1/n4418 ), .C(\MCD/rd_wt_1/n4419 ), .D(\MCD/rd_wt_1/n4420 )
         );
    snl_ao023x1 \MCD/rd_wt_1/U89  ( .Z(ronly1), .A(\stream1[27] ), .B(
        \stream1[26] ), .C(\MCD/rd_wt_1/n4421 ), .D(\MCD/rd_wt_1/n4422 ), .E(
        \MCD/rd_wt_1/n4423 ) );
    snl_and02x1 \MCD/rd_wt_1/U90  ( .Z(po_shelter_h1), .A(\MCD/rd_wt_1/n4424 ), 
        .B(\stream1[25] ) );
    snl_aoi012x1 \MCD/rd_wt_1/U91  ( .ZN(\MCD/rd_wt_1/n4425 ), .A(
        \MCD/rd_wt_1/bacc ), .B(\stream1[1] ), .C(\MCD/rd_wt_1/n4426 ) );
    snl_nor02x1 \MCD/rd_wt_1/U96  ( .ZN(\MCD/rd_wt_1/n4424 ), .A(\stream1[27] 
        ), .B(\stream1[26] ) );
    snl_oai012x1 \MCD/rd_wt_1/U113  ( .ZN(\MCD/rd_wt_1/n4450 ), .A(
        \MCD/rd_wt_1/n4429 ), .B(\MCD/rd_wt_1/n4437 ), .C(\MCD/rd_wt_1/n4451 )
         );
    snl_invx05 \MCD/rd_wt_1/U134  ( .ZN(\MCD/rd_wt_1/n4457 ), .A(
        \MCD/rd_wt_1/n4441 ) );
    snl_invx05 \MCD/rd_wt_1/U98  ( .ZN(\MCD/rd_wt_1/n4438 ), .A(\stream1[26] )
         );
    snl_nor02x1 \MCD/rd_wt_1/U101  ( .ZN(\MCD/rd_wt_1/n4439 ), .A(
        \MCD/rd_wt_1/n4426 ), .B(\stream1[1] ) );
    snl_nand03x0 \MCD/rd_wt_1/U108  ( .ZN(\MCD/rd_wt_1/n4430 ), .A(
        \MCD/rd_wt_1/n4424 ), .B(\MCD/rd_wt_1/n4444 ), .C(\stream1[14] ) );
    snl_nor03x0 \MCD/rd_wt_1/U141  ( .ZN(\MCD/rd_wt_1/n4428 ), .A(
        \MCD/rd_wt_1/n4457 ), .B(\stream1[0] ), .C(\MCD/rd_wt_1/n4443 ) );
    snl_ffqrnx1 \MCD/rd_wt_1/ciff_reg  ( .Q(\MCD/rd_wt_1/ciff ), .D(pk_ciffh), 
        .RN(n10733), .CP(SCLK) );
    snl_nand03x0 \MCD/rd_wt_1/U106  ( .ZN(\MCD/rd_wt_1/n4443 ), .A(
        \stream1[1] ), .B(\MCD/rd_wt_1/n4426 ), .C(\MCD/rd_wt_1/n4432 ) );
    snl_and23x0 \MCD/rd_wt_1/U121  ( .Z(\MCD/rd_wt_1/n4462 ), .A(
        \MCD/rd_wt_1/n4437 ), .B(\stream1[10] ), .C(\MCD/rd_wt_1/n4424 ) );
    snl_nor02x1 \MCD/rd_wt_1/U126  ( .ZN(\MCD/rd_wt_1/n4419 ), .A(ronly1), .B(
        wonly1) );
    snl_nand14x0 \MCD/rd_wt_1/U128  ( .ZN(\MCD/rd_wt_1/n4420 ), .A(
        \stream1[22] ), .B(\MCD/rd_wt_1/n4436 ), .C(\MCD/rd_wt_1/n4423 ), .D(
        \MCD/rd_wt_1/n4450 ) );
    snl_invx05 \MCD/rd_wt_1/U146  ( .ZN(\MCD/rd_wt_1/n4453 ), .A(\stream1[18] 
        ) );
    snl_invx05 \MCD/rd_wt_1/U99  ( .ZN(\MCD/rd_wt_1/n4434 ), .A(
        \MCD/rd_wt_1/bacc ) );
    snl_aoi022x1 \MCD/rd_wt_1/U114  ( .ZN(\MCD/rd_wt_1/n4452 ), .A(
        \MCD/rd_wt_1/n4434 ), .B(\MCD/rd_wt_1/n4453 ), .C(\MCD/rd_wt_1/bacc ), 
        .D(\stream1[18] ) );
    snl_invx05 \MCD/rd_wt_1/U133  ( .ZN(sequencial1), .A(\MCD/rd_wt_1/n4443 )
         );
    snl_invx05 \MCD/rd_wt_1/U107  ( .ZN(\MCD/rd_wt_1/n4444 ), .A(\stream1[15] 
        ) );
    snl_nand02x1 \MCD/rd_wt_1/U120  ( .ZN(\MCD/rd_wt_1/n4460 ), .A(
        \MCD/rd_wt_1/n4443 ), .B(\MCD/rd_wt_1/n4461 ) );
    snl_muxi21x1 \MCD/rd_wt_1/U115  ( .ZN(\MCD/rd_wt_1/n4454 ), .A(
        \MCD/rd_wt_1/n4435 ), .B(\MCD/rd_wt_1/n4425 ), .S(\MCD/rd_wt_1/ciff )
         );
    snl_nor02x1 \MCD/rd_wt_1/U132  ( .ZN(rrmw1), .A(\MCD/rd_wt_1/n4449 ), .B(
        \MCD/rd_wt_1/n4422 ) );
    snl_xor2x0 \MCD/rd_wt_1/U95  ( .Z(\MCD/rd_wt_1/n4436 ), .A(\stream1[21] ), 
        .B(\stream1[20] ) );
    snl_invx05 \MCD/rd_wt_1/U97  ( .ZN(\MCD/rd_wt_1/n4437 ), .A(\stream1[9] )
         );
    snl_invx05 \MCD/rd_wt_1/U109  ( .ZN(\MCD/rd_wt_1/n4445 ), .A(\stream1[13] 
        ) );
    snl_invx05 \MCD/rd_wt_1/U129  ( .ZN(rmw11), .A(\MCD/rd_wt_1/n4420 ) );
    snl_invx05 \MCD/rd_wt_1/U140  ( .ZN(\MCD/rd_wt_1/n4422 ), .A(
        \MCD/rd_wt_1/n4450 ) );
    snl_invx05 \MCD/rd_wt_1/U100  ( .ZN(\MCD/rd_wt_1/n4426 ), .A(\stream1[2] )
         );
    snl_oai113x0 \MCD/rd_wt_1/U112  ( .ZN(\MCD/rd_wt_1/n4449 ), .A(
        \MCD/rd_wt_1/n4441 ), .B(\stream1[0] ), .C(\MCD/rd_wt_1/n4431 ), .D(
        \MCD/rd_wt_1/n4423 ), .E(\MCD/rd_wt_1/n4448 ) );
    snl_invx05 \MCD/rd_wt_1/U135  ( .ZN(\MCD/rd_wt_1/n4435 ), .A(
        \MCD/rd_wt_1/n4439 ) );
    snl_oai013x0 \MCD/rd_wt_1/U110  ( .ZN(\MCD/rd_wt_1/n4423 ), .A(
        \MCD/rd_wt_1/n4444 ), .B(\MCD/rd_wt_1/n4446 ), .C(\MCD/rd_wt_1/n4428 ), 
        .D(\MCD/rd_wt_1/n4447 ) );
    snl_and34x0 \MCD/rd_wt_1/U127  ( .Z(wonly1), .A(\MCD/rd_wt_1/n4423 ), .B(
        \MCD/rd_wt_1/n4422 ), .C(\stream1[22] ), .D(\MCD/rd_wt_1/n4436 ) );
    snl_invx05 \MCD/rd_wt_1/U137  ( .ZN(\MCD/rd_wt_1/n4446 ), .A(
        \MCD/rd_wt_1/n4460 ) );
    snl_invx05 \MCD/rd_wt_1/U102  ( .ZN(\MCD/rd_wt_1/n4440 ), .A(\stream1[0] )
         );
    snl_aoi222x0 \MCD/rd_wt_1/U119  ( .ZN(\MCD/rd_wt_1/n4459 ), .A(
        \MCD/rd_wt_1/n4426 ), .B(\MCD/rd_wt_1/n4442 ), .C(\MCD/rd_wt_1/n4439 ), 
        .D(\MCD/rd_wt_1/n4434 ), .E(\stream1[1] ), .F(\MCD/rd_wt_1/n4441 ) );
    snl_aoi022x1 \MCD/rd_wt_1/U142  ( .ZN(\MCD/rd_wt_1/n4466 ), .A(
        \MCD/rd_wt_1/n4456 ), .B(\MCD/rd_wt_1/n4440 ), .C(\MCD/rd_wt_1/n4455 ), 
        .D(\stream1[0] ) );
    snl_aoi012x1 \MCD/rd_wt_1/U125  ( .ZN(\MCD/rd_wt_1/n4421 ), .A(
        \stream1[19] ), .B(\MCD/rd_wt_1/n4452 ), .C(\stream1[25] ) );
    snl_nor02x1 \MCD/rd_wt_1/U105  ( .ZN(\MCD/rd_wt_1/n4432 ), .A(
        \MCD/rd_wt_1/n4438 ), .B(\stream1[27] ) );
    snl_nor02x1 \MCD/rd_wt_1/U122  ( .ZN(\MCD/rd_wt_1/n4463 ), .A(
        \stream1[13] ), .B(\MCD/rd_wt_1/n4430 ) );
    snl_oa113x1 \MCD/rd_wt_1/U139  ( .Z(\MCD/rd_wt_1/n4429 ), .A(
        \MCD/rd_wt_1/n4465 ), .B(\MCD/rd_wt_1/n4431 ), .C(\MCD/rd_wt_1/n4440 ), 
        .D(\MCD/rd_wt_1/n4443 ), .E(\MCD/rd_wt_1/n4467 ) );
    snl_oa012x1 \MCD/rd_wt_1/U92  ( .Z(\MCD/rd_wt_1/n4427 ), .A(
        \MCD/rd_wt_1/n4428 ), .B(\MCD/rd_wt_1/n4429 ), .C(\MCD/rd_wt_1/n4430 )
         );
    snl_muxi21x1 \MCD/rd_wt_1/U145  ( .ZN(\MCD/rd_wt_1/n4447 ), .A(
        \MCD/rd_wt_1/n4464 ), .B(\MCD/rd_wt_1/n4463 ), .S(\stream1[12] ) );
    snl_nand02x1 \MCD/rd_wt_1/U93  ( .ZN(\MCD/rd_wt_1/n4431 ), .A(
        \MCD/rd_wt_1/n4432 ), .B(\stream1[1] ) );
    snl_invx05 \MCD/rd_wt_1/U104  ( .ZN(\MCD/rd_wt_1/n4442 ), .A(pk_sign_h) );
    snl_aoi222x0 \MCD/rd_wt_1/U117  ( .ZN(\MCD/rd_wt_1/n4456 ), .A(pk_sign_h), 
        .B(\MCD/rd_wt_1/n4426 ), .C(\MCD/rd_wt_1/n4439 ), .D(
        \MCD/rd_wt_1/bacc ), .E(\MCD/rd_wt_1/n4457 ), .F(\stream1[1] ) );
    snl_nand03x0 \MCD/rd_wt_1/U130  ( .ZN(\MCD/rd_wt_1/n4418 ), .A(
        \MCD/rd_wt_1/n4449 ), .B(\MCD/rd_wt_1/n4450 ), .C(\MCD/rd_wt_1/n4448 )
         );
    snl_nand02x1 \MCD/rd_wt_1/U138  ( .ZN(\MCD/rd_wt_1/n4467 ), .A(
        \MCD/rd_wt_1/n4468 ), .B(\MCD/rd_wt_1/n4432 ) );
    snl_aoi013x0 \MCD/rd_wt_1/U116  ( .ZN(\MCD/rd_wt_1/n4455 ), .A(ph_piosl_h), 
        .B(\pk_stat_h[18] ), .C(\stream1[1] ), .D(\MCD/rd_wt_1/n4454 ) );
    snl_nor02x1 \MCD/rd_wt_1/U123  ( .ZN(\MCD/rd_wt_1/n4464 ), .A(
        \MCD/rd_wt_1/n4427 ), .B(\MCD/rd_wt_1/n4445 ) );
    snl_invx05 \MCD/rd_wt_1/U131  ( .ZN(rmw21), .A(\MCD/rd_wt_1/n4418 ) );
    snl_ffqrnx1 \MCD/rd_wt_1/bacc_reg  ( .Q(\MCD/rd_wt_1/bacc ), .D(pk_bacch), 
        .RN(n10733), .CP(SCLK) );
    snl_nor02x1 \MCD/rd_wt_1/U94  ( .ZN(\MCD/rd_wt_1/n4433 ), .A(
        \MCD/rd_wt_1/n4434 ), .B(\MCD/rd_wt_1/n4435 ) );
    snl_aoi022x1 \MCD/rd_wt_1/U143  ( .ZN(\MCD/rd_wt_1/n4468 ), .A(
        \MCD/rd_wt_1/n4459 ), .B(\MCD/rd_wt_1/n4440 ), .C(\MCD/rd_wt_1/n4458 ), 
        .D(\stream1[0] ) );
    snl_muxi21x1 \MCD/rd_wt_1/U144  ( .ZN(\MCD/rd_wt_1/n4451 ), .A(
        \MCD/rd_wt_1/n4462 ), .B(\MCD/rd_wt_1/n4460 ), .S(\stream1[11] ) );
    snl_nand12x1 \MCD/rd_wt_1/U103  ( .ZN(\MCD/rd_wt_1/n4441 ), .A(pk_pcon31_h
        ), .B(\MCD/rd_wt_1/ciff ) );
    snl_nor03x0 \MCD/rd_wt_1/U111  ( .ZN(\MCD/rd_wt_1/n4448 ), .A(
        \stream1[22] ), .B(\stream1[20] ), .C(\stream1[21] ) );
    snl_nand02x1 \MCD/rd_wt_1/U136  ( .ZN(\MCD/rd_wt_1/n4461 ), .A(
        \MCD/rd_wt_1/n4466 ), .B(\MCD/rd_wt_1/n4432 ) );
    snl_ao022x1 \MCD/rd_wt_1/U124  ( .Z(\MCD/rd_wt_1/n4465 ), .A(
        \MCD/rd_wt_1/bacc ), .B(\MCD/rd_wt_1/ciff ), .C(\pk_stat_h[18] ), .D(
        ph_piosl_h) );
    snl_muxi21x1 \MCD/rd_wt_1/U118  ( .ZN(\MCD/rd_wt_1/n4458 ), .A(
        \MCD/rd_wt_1/n4426 ), .B(\MCD/rd_wt_1/n4433 ), .S(\MCD/rd_wt_1/ciff )
         );
    snl_mux21x1 \ADOSEL/seladr_4/U10  ( .Z(LOUT[31]), .A(1'b0), .B(
        \pgmuxout[31] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U12  ( .Z(LOUT[29]), .A(1'b1), .B(
        \pgmuxout[29] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U13  ( .Z(LOUT[28]), .A(1'b0), .B(
        \pgmuxout[28] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U14  ( .Z(LOUT[27]), .A(\pgsadrh[27] ), .B(
        \pgmuxout[27] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U15  ( .Z(LOUT[26]), .A(\pgsadrh[26] ), .B(
        \pgmuxout[26] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U17  ( .Z(LOUT[24]), .A(\pgsadrh[24] ), .B(
        \pgmuxout[24] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U11  ( .Z(LOUT[30]), .A(1'b1), .B(
        \pgmuxout[30] ), .S(ph_ldaoutenh4) );
    snl_mux21x1 \ADOSEL/seladr_4/U16  ( .Z(LOUT[25]), .A(\pgsadrh[25] ), .B(
        \pgmuxout[25] ), .S(ph_ldaoutenh4) );
    snl_nand12x1 \MAIN/STM/U14  ( .ZN(\MAIN/STM/exestage_err ), .A(
        \MAIN/ADROVH ), .B(\MAIN/STM/n3365 ) );
    snl_nor02x1 \MAIN/STM/U13  ( .ZN(pgbnolth), .A(stage_2), .B(
        \MAIN/STM/n3366 ) );
    snl_nor02x1 \MAIN/STM/U12  ( .ZN(\MAIN/STM/n3365 ), .A(\MAIN/STM/exe_err3 
        ), .B(\MAIN/STM/exe_err2 ) );
    snl_nand02x1 \MAIN/STM/U10  ( .ZN(lbus_start), .A(\MAIN/STM/sa_start2 ), 
        .B(\MAIN/STM/sa_start3 ) );
    snl_nand12x1 \MAIN/STM/U15  ( .ZN(ph_filewr_h), .A(
        \MAIN/STM/srgfilewren_h ), .B(\MAIN/STM/n3364 ) );
    snl_nor03x0 \MAIN/STM/U17  ( .ZN(\MAIN/STM/n3364 ), .A(
        \MAIN/STM/exec_eoc3 ), .B(\MAIN/STM/exec_eoc2 ), .C(
        \MAIN/STM/exec_eoc1 ) );
    snl_nand12x1 \MAIN/STM/U11  ( .ZN(\MAIN/exe_end ), .A(\MAIN/STM/exec_eoc ), 
        .B(\MAIN/STM/n3364 ) );
    snl_invx05 \MAIN/STM/U19  ( .ZN(\MAIN/STM/execute_err ), .A(
        \MAIN/STM/n3365 ) );
    snl_or03x1 \MAIN/STM/U16  ( .Z(\MAIN/STM/seq_end ), .A(
        \MAIN/STM/exec_end1 ), .B(\MAIN/STM/exec_end2 ), .C(
        \MAIN/STM/exec_end3 ) );
    snl_invx05 \MAIN/STM/U18  ( .ZN(\MAIN/STM/n3366 ), .A(\MAIN/STM/bnolth )
         );
    snl_nand12x1 \MAIN/SW/U29  ( .ZN(\MAIN/SW/nst[0] ), .A(polcore_end), .B(
        \MAIN/SW/n3322 ) );
    snl_ffqrnx1 \MAIN/SW/wst_reg[0]  ( .Q(\MAIN/SW/wst[0] ), .D(
        \MAIN/SW/nst[0] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \MAIN/SW/U30  ( .ZN(\MAIN/SW/n3323 ), .A(\MAIN/SW/wst[0] ) );
    snl_nand02x1 \MAIN/SW/U32  ( .ZN(\MAIN/SW/n3322 ), .A(\MAIN/st_swctl ), 
        .B(\MAIN/SW/n3323 ) );
    snl_ffqrnx1 \MAIN/SW/wst_reg[1]  ( .Q(\MAIN/sw_end ), .D(polcore_end), 
        .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nor02x1 \MAIN/SW/U31  ( .ZN(polcore_end), .A(\MAIN/SW/n3323 ), .B(
        \MAIN/sw_end ) );
    snl_ffqx1 \MAIN/SW/excep_enable_reg  ( .Q(\MAIN/excep_enable ), .D(
        \MAIN/SW/nst[0] ), .CP(SCLK) );
    snl_mux21x1 \ADOSEL/seladr_3/U10  ( .Z(LOUT[23]), .A(\pgsadrh[23] ), .B(
        \pgmuxout[23] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U12  ( .Z(LOUT[21]), .A(\pgsadrh[21] ), .B(
        \pgmuxout[21] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U13  ( .Z(LOUT[20]), .A(\pgsadrh[20] ), .B(
        \pgmuxout[20] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U14  ( .Z(LOUT[19]), .A(\pgsadrh[19] ), .B(
        \pgmuxout[19] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U15  ( .Z(LOUT[18]), .A(\pgsadrh[18] ), .B(
        \pgmuxout[18] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U17  ( .Z(LOUT[16]), .A(\pgsadrh[16] ), .B(
        \pgmuxout[16] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U11  ( .Z(LOUT[22]), .A(\pgsadrh[22] ), .B(
        \pgmuxout[22] ), .S(ph_ldaoutenh3) );
    snl_mux21x1 \ADOSEL/seladr_3/U16  ( .Z(LOUT[17]), .A(\pgsadrh[17] ), .B(
        \pgmuxout[17] ), .S(ph_ldaoutenh3) );
    snl_bufx2 \CODEQ/phque12_1/U265  ( .Z(\CODEQ/phque12_1/n767 ), .A(n10731)
         );
    snl_or02x1 \CODEQ/phque12_1/U271  ( .Z(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .A(step3_cf), .B(step1_cf)
         );
    snl_invx05 \CODEQ/phque12_1/U338  ( .ZN(\CODEQ/nqueue1[35] ), .A(
        \CODEQ/phque12_1/queue1[35] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[31]  ( .Q(
        \CODEQ/phque12_1/queue1[31] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[31]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[28]  ( .Q(
        \CODEQ/phque12_1/queue1[28] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[28]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U356  ( .ZN(\CODEQ/nqueue1[55] ), .A(
        \CODEQ/phque12_1/queue1[55] ) );
    snl_invx05 \CODEQ/phque12_1/U371  ( .ZN(\CODEQ/nqueue2[1] ), .A(
        \CODEQ/phque12_1/queue2[1] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[30]  ( .Q(
        \CODEQ/phque12_1/queue2[30] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[30]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[29]  ( .Q(
        \CODEQ/phque12_1/queue2[29] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[29]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U276  ( .ZN(\CODEQ/nqueue1[27] ), .A(
        \CODEQ/phque12_1/queue1[27] ) );
    snl_invx05 \CODEQ/phque12_1/U278  ( .ZN(\CODEQ/nqueue2[40] ), .A(
        \CODEQ/phque12_1/queue2[40] ) );
    snl_invx05 \CODEQ/phque12_1/U286  ( .ZN(\CODEQ/nqueue2[37] ), .A(
        \CODEQ/phque12_1/queue2[37] ) );
    snl_invx05 \CODEQ/phque12_1/U294  ( .ZN(\CODEQ/nqueue1[47] ), .A(
        \stream1[15] ) );
    snl_invx05 \CODEQ/phque12_1/U304  ( .ZN(\CODEQ/nqueue2[24] ), .A(
        \CODEQ/phque12_1/queue2[24] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[12]  ( .Q(
        \CODEQ/phque12_1/queue1[12] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[12]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[39]  ( .Q(
        \CODEQ/phque12_1/queue2[39] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[39]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[13]  ( .Q(
        \CODEQ/phque12_1/queue2[13] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[13]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[20]  ( .Q(
        \CODEQ/phque12_1/queue2[20] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[20]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[6]  ( .Q(
        \CODEQ/phque12_1/queue2[6] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[6]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U323  ( .ZN(\CODEQ/nqueue2[27] ), .A(
        \CODEQ/phque12_1/queue2[27] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[38]  ( .Q(
        \CODEQ/phque12_1/queue1[38] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[38]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[21]  ( .Q(
        \CODEQ/phque12_1/queue1[21] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[21]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[34]  ( .Q(\stream2[2] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[34]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U316  ( .ZN(\CODEQ/nqueue1[53] ), .A(
        \stream1[21] ) );
    snl_invx05 \CODEQ/phque12_1/U331  ( .ZN(\CODEQ/nqueue1[45] ), .A(
        \stream1[13] ) );
    snl_invx05 \CODEQ/phque12_1/U378  ( .ZN(\CODEQ/nqueue2[16] ), .A(
        \CODEQ/phque12_1/queue2[16] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[35]  ( .Q(
        \CODEQ/phque12_1/queue1[35] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[35]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U281  ( .ZN(\CODEQ/nqueue2[11] ), .A(
        \CODEQ/phque12_1/queue2[11] ) );
    snl_invx05 \CODEQ/phque12_1/U311  ( .ZN(\CODEQ/nqueue2[12] ), .A(
        \CODEQ/phque12_1/queue2[12] ) );
    snl_invx05 \CODEQ/phque12_1/U336  ( .ZN(\CODEQ/nqueue2[31] ), .A(
        \CODEQ/phque12_1/queue2[31] ) );
    snl_invx05 \CODEQ/phque12_1/U343  ( .ZN(\CODEQ/nqueue2[2] ), .A(
        \CODEQ/phque12_1/queue2[2] ) );
    snl_invx05 \CODEQ/phque12_1/U344  ( .ZN(\CODEQ/nqueue2[29] ), .A(
        \CODEQ/phque12_1/queue2[29] ) );
    snl_invx05 \CODEQ/phque12_1/U363  ( .ZN(\CODEQ/nqueue1[49] ), .A(
        \CODEQ/phque12_1/queue1[49] ) );
    snl_invx05 \CODEQ/phque12_1/U381  ( .ZN(\CODEQ/nqueue1[29] ), .A(
        \CODEQ/phque12_1/queue1[29] ) );
    snl_invx05 \CODEQ/phque12_1/U386  ( .ZN(\CODEQ/nqueue2[54] ), .A(
        \stream2[22] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[25]  ( .Q(
        \CODEQ/phque12_1/queue1[25] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[25]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[16]  ( .Q(
        \CODEQ/phque12_1/queue1[16] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[16]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[24]  ( .Q(
        \CODEQ/phque12_1/queue2[24] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[24]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[17]  ( .Q(
        \CODEQ/phque12_1/queue2[17] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[17]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[2]  ( .Q(
        \CODEQ/phque12_1/queue2[2] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[2]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[26]  ( .Q(
        \CODEQ/phque12_1/queue2[26] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[26]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[15]  ( .Q(
        \CODEQ/phque12_1/queue2[15] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[15]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[0]  ( .Q(
        \CODEQ/phque12_1/queue2[0] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[0]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U358  ( .ZN(\CODEQ/nqueue1[8] ), .A(
        \CODEQ/phque12_1/queue1[8] ) );
    snl_invx05 \CODEQ/phque12_1/U364  ( .ZN(\CODEQ/nqueue2[8] ), .A(
        \CODEQ/phque12_1/queue2[8] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[14]  ( .Q(
        \CODEQ/phque12_1/queue1[14] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[14]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[27]  ( .Q(
        \CODEQ/phque12_1/queue1[27] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[27]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[37]  ( .Q(
        \CODEQ/phque12_1/queue1[37] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[37]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[36]  ( .Q(
        \CODEQ/phque12_1/queue2[36] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[36]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[9]  ( .Q(
        \CODEQ/phque12_1/queue2[9] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[9]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U293  ( .ZN(\CODEQ/nqueue1[50] ), .A(
        \stream1[18] ) );
    snl_invx05 \CODEQ/phque12_1/U324  ( .ZN(\CODEQ/nqueue2[36] ), .A(
        \CODEQ/phque12_1/queue2[36] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[23]  ( .Q(
        \CODEQ/phque12_1/queue1[23] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[23]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[10]  ( .Q(
        \CODEQ/phque12_1/queue1[10] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[10]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U303  ( .ZN(\CODEQ/nqueue2[7] ), .A(
        \CODEQ/phque12_1/queue2[7] ) );
    snl_invx05 \CODEQ/phque12_1/U388  ( .ZN(\CODEQ/nqueue2[28] ), .A(
        \CODEQ/phque12_1/queue2[28] ) );
    snl_invx05 \CODEQ/phque12_1/U280  ( .ZN(\CODEQ/nqueue1[59] ), .A(
        \stream1[27] ) );
    snl_invx05 \CODEQ/phque12_1/U288  ( .ZN(\CODEQ/nqueue2[25] ), .A(
        \CODEQ/phque12_1/queue2[25] ) );
    snl_invx05 \CODEQ/phque12_1/U351  ( .ZN(\CODEQ/nqueue1[15] ), .A(
        \CODEQ/phque12_1/queue1[15] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[22]  ( .Q(
        \CODEQ/phque12_1/queue2[22] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[22]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[11]  ( .Q(
        \CODEQ/phque12_1/queue2[11] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[11]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[4]  ( .Q(
        \CODEQ/phque12_1/queue2[4] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[4]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U376  ( .ZN(\CODEQ/nqueue2[30] ), .A(
        \CODEQ/phque12_1/queue2[30] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[33]  ( .Q(\stream1[1] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[33]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[32]  ( .Q(\stream2[0] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[32]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[18]  ( .Q(
        \CODEQ/phque12_1/queue2[18] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[18]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[19]  ( .Q(
        \CODEQ/phque12_1/queue1[19] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[19]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U318  ( .ZN(\CODEQ/nqueue2[19] ), .A(
        \CODEQ/phque12_1/queue2[19] ) );
    snl_invx05 \CODEQ/phque12_1/U337  ( .ZN(\CODEQ/nqueue1[28] ), .A(
        \CODEQ/phque12_1/queue1[28] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[57]  ( .Q(\stream2[25] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[57]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U310  ( .ZN(\CODEQ/nqueue1[6] ), .A(
        \CODEQ/phque12_1/queue1[6] ) );
    snl_invx05 \CODEQ/phque12_1/U359  ( .ZN(\CODEQ/nqueue1[23] ), .A(
        \CODEQ/phque12_1/queue1[23] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[7]  ( .Q(
        \CODEQ/phque12_1/queue1[7] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[7]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[56]  ( .Q(
        \CODEQ/phque12_1/queue1[56] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[56]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_bufx2 \CODEQ/phque12_1/U266  ( .Z(\CODEQ/phque12_1/n769 ), .A(n10731)
         );
    snl_bufx2 \CODEQ/phque12_1/U267  ( .Z(\CODEQ/phque12_1/n768 ), .A(n10731)
         );
    snl_or02x1 \CODEQ/phque12_1/U269  ( .Z(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .A(step4_cf), .B(step2_cf)
         );
    snl_bufx1 \CODEQ/phque12_1/U270  ( .Z(\CODEQ/phque12_1/n771 ), .A(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ) );
    snl_invx05 \CODEQ/phque12_1/U277  ( .ZN(\CODEQ/nqueue1[32] ), .A(
        \stream1[0] ) );
    snl_invx05 \CODEQ/phque12_1/U289  ( .ZN(\CODEQ/nqueue2[34] ), .A(
        \stream2[2] ) );
    snl_invx05 \CODEQ/phque12_1/U319  ( .ZN(\CODEQ/nqueue2[48] ), .A(
        \CODEQ/phque12_1/queue2[48] ) );
    snl_invx05 \CODEQ/phque12_1/U342  ( .ZN(\CODEQ/nqueue2[55] ), .A(
        \CODEQ/phque12_1/queue2[55] ) );
    snl_invx05 \CODEQ/phque12_1/U365  ( .ZN(\CODEQ/nqueue2[23] ), .A(
        \CODEQ/phque12_1/queue2[23] ) );
    snl_invx05 \CODEQ/phque12_1/U380  ( .ZN(\CODEQ/nqueue1[2] ), .A(
        \CODEQ/phque12_1/queue1[2] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[46]  ( .Q(\stream1[14] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[46]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[47]  ( .Q(\stream2[15] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[47]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[52]  ( .Q(\stream1[20] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[52]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U350  ( .ZN(\CODEQ/nqueue1[1] ), .A(
        \CODEQ/phque12_1/queue1[1] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[3]  ( .Q(
        \CODEQ/phque12_1/queue1[3] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[3]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U377  ( .ZN(\CODEQ/nqueue1[54] ), .A(
        \stream1[22] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[53]  ( .Q(\stream2[21] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[53]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U292  ( .ZN(\CODEQ/nqueue1[30] ), .A(
        \CODEQ/phque12_1/queue1[30] ) );
    snl_invx05 \CODEQ/phque12_1/U302  ( .ZN(\CODEQ/nqueue1[46] ), .A(
        \stream1[14] ) );
    snl_invx05 \CODEQ/phque12_1/U325  ( .ZN(\CODEQ/nqueue2[53] ), .A(
        \stream2[21] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[43]  ( .Q(\stream2[11] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[43]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[42]  ( .Q(\stream1[10] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[42]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U295  ( .ZN(\CODEQ/nqueue2[50] ), .A(
        \stream2[18] ) );
    snl_invx05 \CODEQ/phque12_1/U389  ( .ZN(\CODEQ/nqueue1[17] ), .A(
        \CODEQ/phque12_1/queue1[17] ) );
    snl_invx05 \CODEQ/phque12_1/U305  ( .ZN(\CODEQ/nqueue2[58] ), .A(
        \stream2[26] ) );
    snl_invx05 \CODEQ/phque12_1/U322  ( .ZN(\CODEQ/nqueue2[4] ), .A(
        \CODEQ/phque12_1/queue2[4] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[59]  ( .Q(\stream1[27] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[59]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[40]  ( .Q(
        \CODEQ/phque12_1/queue1[40] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[40]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[8]  ( .Q(
        \CODEQ/phque12_1/queue1[8] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[8]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U279  ( .ZN(\CODEQ/nqueue1[44] ), .A(
        \stream1[12] ) );
    snl_invx05 \CODEQ/phque12_1/U339  ( .ZN(\CODEQ/nqueue1[21] ), .A(
        \CODEQ/phque12_1/queue1[21] ) );
    snl_invx05 \CODEQ/phque12_1/U357  ( .ZN(\CODEQ/nqueue2[14] ), .A(
        \CODEQ/phque12_1/queue2[14] ) );
    snl_invx05 \CODEQ/phque12_1/U370  ( .ZN(\CODEQ/nqueue2[44] ), .A(
        \stream2[12] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[58]  ( .Q(\stream2[26] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[58]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[41]  ( .Q(\stream2[9] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[41]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[50]  ( .Q(\stream1[18] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[50]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[51]  ( .Q(\stream2[19] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[51]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[48]  ( .Q(
        \CODEQ/phque12_1/queue2[48] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[48]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[49]  ( .Q(
        \CODEQ/phque12_1/queue1[49] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[49]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U387  ( .ZN(\CODEQ/nqueue2[3] ), .A(
        \CODEQ/phque12_1/queue2[3] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[1]  ( .Q(
        \CODEQ/phque12_1/queue1[1] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[1]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[45]  ( .Q(\stream2[13] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[45]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U287  ( .ZN(\CODEQ/nqueue2[6] ), .A(
        \CODEQ/phque12_1/queue2[6] ) );
    snl_invx05 \CODEQ/phque12_1/U317  ( .ZN(\CODEQ/nqueue1[11] ), .A(
        \CODEQ/phque12_1/queue1[11] ) );
    snl_invx05 \CODEQ/phque12_1/U345  ( .ZN(\CODEQ/nqueue2[33] ), .A(
        \stream2[1] ) );
    snl_invx05 \CODEQ/phque12_1/U362  ( .ZN(\CODEQ/nqueue1[0] ), .A(
        \CODEQ/phque12_1/queue1[0] ) );
    snl_invx05 \CODEQ/phque12_1/U379  ( .ZN(\CODEQ/nqueue2[21] ), .A(
        \CODEQ/phque12_1/queue2[21] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[44]  ( .Q(\stream1[12] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[44]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[5]  ( .Q(
        \CODEQ/phque12_1/queue1[5] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[5]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[54]  ( .Q(\stream1[22] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[54]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[55]  ( .Q(
        \CODEQ/phque12_1/queue2[55] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[55]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U330  ( .ZN(\CODEQ/nqueue2[41] ), .A(
        \stream2[9] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[44]  ( .Q(\stream2[12] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[44]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U272  ( .ZN(\CODEQ/nqueue2[49] ), .A(
        \CODEQ/phque12_1/queue2[49] ) );
    snl_invx05 \CODEQ/phque12_1/U355  ( .ZN(\CODEQ/nqueue2[0] ), .A(
        \CODEQ/phque12_1/queue2[0] ) );
    snl_invx05 \CODEQ/phque12_1/U369  ( .ZN(\CODEQ/nqueue2[15] ), .A(
        \CODEQ/phque12_1/queue2[15] ) );
    snl_invx05 \CODEQ/phque12_1/U372  ( .ZN(\CODEQ/nqueue1[9] ), .A(
        \CODEQ/phque12_1/queue1[9] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[45]  ( .Q(\stream1[13] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[45]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[4]  ( .Q(
        \CODEQ/phque12_1/queue1[4] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[4]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U285  ( .ZN(\CODEQ/nqueue1[19] ), .A(
        \CODEQ/phque12_1/queue1[19] ) );
    snl_invx05 \CODEQ/phque12_1/U297  ( .ZN(\CODEQ/nqueue1[52] ), .A(
        \stream1[20] ) );
    snl_invx05 \CODEQ/phque12_1/U320  ( .ZN(\CODEQ/nqueue1[5] ), .A(
        \CODEQ/phque12_1/queue1[5] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[55]  ( .Q(
        \CODEQ/phque12_1/queue1[55] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[55]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[54]  ( .Q(\stream2[22] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[54]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U307  ( .ZN(\CODEQ/nqueue2[35] ), .A(
        \CODEQ/phque12_1/queue2[35] ) );
    snl_invx05 \CODEQ/phque12_1/U315  ( .ZN(\CODEQ/nqueue1[38] ), .A(
        \CODEQ/phque12_1/queue1[38] ) );
    snl_invx05 \CODEQ/phque12_1/U332  ( .ZN(\CODEQ/nqueue2[17] ), .A(
        \CODEQ/phque12_1/queue2[17] ) );
    snl_invx05 \CODEQ/phque12_1/U299  ( .ZN(\CODEQ/nqueue2[13] ), .A(
        \CODEQ/phque12_1/queue2[13] ) );
    snl_invx05 \CODEQ/phque12_1/U329  ( .ZN(\CODEQ/nqueue2[10] ), .A(
        \CODEQ/phque12_1/queue2[10] ) );
    snl_invx05 \CODEQ/phque12_1/U347  ( .ZN(\CODEQ/nqueue2[9] ), .A(
        \CODEQ/phque12_1/queue2[9] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[58]  ( .Q(\stream1[26] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[58]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[41]  ( .Q(\stream1[9] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[41]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[9]  ( .Q(
        \CODEQ/phque12_1/queue1[9] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[9]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[59]  ( .Q(\stream2[27] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[59]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[40]  ( .Q(
        \CODEQ/phque12_1/queue2[40] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[40]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U360  ( .ZN(\CODEQ/nqueue2[45] ), .A(
        \stream2[13] ) );
    snl_invx05 \CODEQ/phque12_1/U385  ( .ZN(\CODEQ/nqueue2[47] ), .A(
        \stream2[15] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[51]  ( .Q(\stream1[19] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[51]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[48]  ( .Q(
        \CODEQ/phque12_1/queue1[48] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[48]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[50]  ( .Q(\stream2[18] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[50]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[49]  ( .Q(
        \CODEQ/phque12_1/queue2[49] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[49]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[0]  ( .Q(
        \CODEQ/phque12_1/queue1[0] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[0]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U382  ( .ZN(\CODEQ/nqueue1[34] ), .A(
        \stream1[2] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[53]  ( .Q(\stream1[21] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[53]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[2]  ( .Q(
        \CODEQ/phque12_1/queue1[2] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[2]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U309  ( .ZN(\CODEQ/nqueue1[31] ), .A(
        \CODEQ/phque12_1/queue1[31] ) );
    snl_invx05 \CODEQ/phque12_1/U340  ( .ZN(\CODEQ/nqueue1[43] ), .A(
        \stream1[11] ) );
    snl_invx05 \CODEQ/phque12_1/U367  ( .ZN(\CODEQ/nqueue2[57] ), .A(
        \stream2[25] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[52]  ( .Q(\stream2[20] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[52]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U275  ( .ZN(\CODEQ/nqueue1[10] ), .A(
        \CODEQ/phque12_1/queue1[10] ) );
    snl_invx05 \CODEQ/phque12_1/U282  ( .ZN(\CODEQ/nqueue2[5] ), .A(
        \CODEQ/phque12_1/queue2[5] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[42]  ( .Q(\stream2[10] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[42]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U290  ( .ZN(\CODEQ/nqueue2[59] ), .A(
        \stream2[27] ) );
    snl_invx05 \CODEQ/phque12_1/U300  ( .ZN(\CODEQ/nqueue2[42] ), .A(
        \stream2[10] ) );
    snl_invx05 \CODEQ/phque12_1/U312  ( .ZN(\CODEQ/nqueue2[51] ), .A(
        \stream2[19] ) );
    snl_invx05 \CODEQ/phque12_1/U335  ( .ZN(\CODEQ/nqueue2[20] ), .A(
        \CODEQ/phque12_1/queue2[20] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[43]  ( .Q(\stream1[11] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[43]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[56]  ( .Q(
        \CODEQ/phque12_1/queue2[56] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[56]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U327  ( .ZN(\CODEQ/nqueue1[51] ), .A(
        \stream1[19] ) );
    snl_invx05 \CODEQ/phque12_1/U349  ( .ZN(\CODEQ/nqueue2[56] ), .A(
        \CODEQ/phque12_1/queue2[56] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[57]  ( .Q(\stream1[25] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[57]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[6]  ( .Q(
        \CODEQ/phque12_1/queue1[6] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[6]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U283  ( .ZN(\CODEQ/nqueue2[26] ), .A(
        \CODEQ/phque12_1/queue2[26] ) );
    snl_invx05 \CODEQ/phque12_1/U313  ( .ZN(\CODEQ/nqueue1[25] ), .A(
        \CODEQ/phque12_1/queue1[25] ) );
    snl_invx05 \CODEQ/phque12_1/U352  ( .ZN(\CODEQ/nqueue1[16] ), .A(
        \CODEQ/phque12_1/queue1[16] ) );
    snl_invx05 \CODEQ/phque12_1/U375  ( .ZN(\CODEQ/nqueue1[40] ), .A(
        \CODEQ/phque12_1/queue1[40] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[47]  ( .Q(\stream1[15] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[47]), .SE(
        \CODEQ/phque12_1/n771 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U390  ( .ZN(\CODEQ/nqueue1[20] ), .A(
        \CODEQ/phque12_1/queue1[20] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[46]  ( .Q(\stream2[14] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n768 ), .SD(CDIN[46]), .SE(
        \CODEQ/phque12_1/n770 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U334  ( .ZN(\CODEQ/nqueue1[3] ), .A(
        \CODEQ/phque12_1/queue1[3] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[11]  ( .Q(
        \CODEQ/phque12_1/queue1[11] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[11]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[22]  ( .Q(
        \CODEQ/phque12_1/queue1[22] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[22]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_bufx1 \CODEQ/phque12_1/U268  ( .Z(\CODEQ/phque12_1/n770 ), .A(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ) );
    snl_invx05 \CODEQ/phque12_1/U273  ( .ZN(\CODEQ/nqueue2[18] ), .A(
        \CODEQ/phque12_1/queue2[18] ) );
    snl_invx05 \CODEQ/phque12_1/U274  ( .ZN(\CODEQ/nqueue1[4] ), .A(
        \CODEQ/phque12_1/queue1[4] ) );
    snl_invx05 \CODEQ/phque12_1/U298  ( .ZN(\CODEQ/nqueue1[7] ), .A(
        \CODEQ/phque12_1/queue1[7] ) );
    snl_invx05 \CODEQ/phque12_1/U308  ( .ZN(\CODEQ/nqueue2[43] ), .A(
        \stream2[11] ) );
    snl_invx05 \CODEQ/phque12_1/U341  ( .ZN(\CODEQ/nqueue1[56] ), .A(
        \CODEQ/phque12_1/queue1[56] ) );
    snl_invx05 \CODEQ/phque12_1/U366  ( .ZN(\CODEQ/nqueue2[32] ), .A(
        \stream2[0] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[23]  ( .Q(
        \CODEQ/phque12_1/queue2[23] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[23]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[10]  ( .Q(
        \CODEQ/phque12_1/queue2[10] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[10]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[5]  ( .Q(
        \CODEQ/phque12_1/queue2[5] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[5]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U383  ( .ZN(\CODEQ/nqueue1[57] ), .A(
        \stream1[25] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[32]  ( .Q(\stream1[0] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n769 ), .SD(CDIN[32]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[33]  ( .Q(\stream2[1] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[33]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[19]  ( .Q(
        \CODEQ/phque12_1/queue2[19] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[19]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[18]  ( .Q(
        \CODEQ/phque12_1/queue1[18] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[18]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U348  ( .ZN(\CODEQ/nqueue2[22] ), .A(
        \CODEQ/phque12_1/queue2[22] ) );
    snl_invx05 \CODEQ/phque12_1/U353  ( .ZN(\CODEQ/nqueue1[36] ), .A(
        \CODEQ/phque12_1/queue1[36] ) );
    snl_invx05 \CODEQ/phque12_1/U374  ( .ZN(\CODEQ/nqueue1[37] ), .A(
        \CODEQ/phque12_1/queue1[37] ) );
    snl_invx05 \CODEQ/phque12_1/U391  ( .ZN(\CODEQ/nqueue1[42] ), .A(
        \stream1[10] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[27]  ( .Q(
        \CODEQ/phque12_1/queue2[27] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[27]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[14]  ( .Q(
        \CODEQ/phque12_1/queue2[14] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[14]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[1]  ( .Q(
        \CODEQ/phque12_1/queue2[1] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[1]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[26]  ( .Q(
        \CODEQ/phque12_1/queue1[26] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[26]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[15]  ( .Q(
        \CODEQ/phque12_1/queue1[15] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[15]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[36]  ( .Q(
        \CODEQ/phque12_1/queue1[36] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[36]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U291  ( .ZN(\CODEQ/nqueue1[12] ), .A(
        \CODEQ/phque12_1/queue1[12] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[37]  ( .Q(
        \CODEQ/phque12_1/queue2[37] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[37]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[8]  ( .Q(
        \CODEQ/phque12_1/queue2[8] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[8]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U296  ( .ZN(\CODEQ/nqueue1[39] ), .A(
        \CODEQ/phque12_1/queue1[39] ) );
    snl_invx05 \CODEQ/phque12_1/U301  ( .ZN(\CODEQ/nqueue1[24] ), .A(
        \CODEQ/phque12_1/queue1[24] ) );
    snl_invx05 \CODEQ/phque12_1/U306  ( .ZN(\CODEQ/nqueue1[13] ), .A(
        \CODEQ/phque12_1/queue1[13] ) );
    snl_invx05 \CODEQ/phque12_1/U321  ( .ZN(\CODEQ/nqueue1[26] ), .A(
        \CODEQ/phque12_1/queue1[26] ) );
    snl_invx05 \CODEQ/phque12_1/U326  ( .ZN(\CODEQ/nqueue1[18] ), .A(
        \CODEQ/phque12_1/queue1[18] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[35]  ( .Q(
        \CODEQ/phque12_1/queue2[35] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[35]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U368  ( .ZN(\CODEQ/nqueue1[14] ), .A(
        \CODEQ/phque12_1/queue1[14] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[34]  ( .Q(\stream1[2] ), .D(
        1'b0), .EN(1'b1), .RN(\CODEQ/phque12_1/n767 ), .SD(CDIN[34]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U284  ( .ZN(\CODEQ/nqueue2[52] ), .A(
        \stream2[20] ) );
    snl_invx05 \CODEQ/phque12_1/U328  ( .ZN(\CODEQ/nqueue1[58] ), .A(
        \stream1[26] ) );
    snl_invx05 \CODEQ/phque12_1/U354  ( .ZN(\CODEQ/nqueue1[48] ), .A(
        \CODEQ/phque12_1/queue1[48] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[17]  ( .Q(
        \CODEQ/phque12_1/queue1[17] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[17]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U373  ( .ZN(\CODEQ/nqueue1[22] ), .A(
        \CODEQ/phque12_1/queue1[22] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[24]  ( .Q(
        \CODEQ/phque12_1/queue1[24] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[24]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U384  ( .ZN(\CODEQ/nqueue2[39] ), .A(
        \CODEQ/phque12_1/queue2[39] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[30]  ( .Q(
        \CODEQ/phque12_1/queue1[30] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[30]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[29]  ( .Q(
        \CODEQ/phque12_1/queue1[29] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[29]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[25]  ( .Q(
        \CODEQ/phque12_1/queue2[25] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[25]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[16]  ( .Q(
        \CODEQ/phque12_1/queue2[16] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[16]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[3]  ( .Q(
        \CODEQ/phque12_1/queue2[3] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[3]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U333  ( .ZN(\CODEQ/nqueue2[46] ), .A(
        \stream2[14] ) );
    snl_invx05 \CODEQ/phque12_1/U346  ( .ZN(\CODEQ/nqueue2[38] ), .A(
        \CODEQ/phque12_1/queue2[38] ) );
    snl_invx05 \CODEQ/phque12_1/U361  ( .ZN(\CODEQ/nqueue1[41] ), .A(
        \stream1[9] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[38]  ( .Q(
        \CODEQ/phque12_1/queue2[38] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[38]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[31]  ( .Q(
        \CODEQ/phque12_1/queue2[31] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[31]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[28]  ( .Q(
        \CODEQ/phque12_1/queue2[28] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[28]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[21]  ( .Q(
        \CODEQ/phque12_1/queue2[21] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[21]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[12]  ( .Q(
        \CODEQ/phque12_1/queue2[12] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[12]), .SE(\CODEQ/phque12_1/n770 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue2_reg[7]  ( .Q(
        \CODEQ/phque12_1/queue2[7] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n768 ), .SD(CDIN[7]), .SE(
        \CODEQ/phque12_1/*cell*3975/U2/CONTROL1 ), .CP(SCLK) );
    snl_invx05 \CODEQ/phque12_1/U314  ( .ZN(\CODEQ/nqueue1[33] ), .A(
        \stream1[1] ) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[39]  ( .Q(
        \CODEQ/phque12_1/queue1[39] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[39]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[20]  ( .Q(
        \CODEQ/phque12_1/queue1[20] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n769 ), .SD(CDIN[20]), .SE(\CODEQ/phque12_1/n771 ), 
        .CP(SCLK) );
    snl_sffqenrnx1 \CODEQ/phque12_1/queue1_reg[13]  ( .Q(
        \CODEQ/phque12_1/queue1[13] ), .D(1'b0), .EN(1'b1), .RN(
        \CODEQ/phque12_1/n767 ), .SD(CDIN[13]), .SE(
        \CODEQ/phque12_1/*cell*3975/U1/CONTROL1 ), .CP(SCLK) );
    snl_invx1 \SADR/SELSEG/U10  ( .ZN(\SADR/SELSEG/n9104 ), .A(
        \SADR/SELSEG/n9084 ) );
    snl_invx1 \SADR/SELSEG/U12  ( .ZN(\SADR/SELSEG/n9099 ), .A(
        \SADR/SELSEG/n9076 ) );
    snl_invx1 \SADR/SELSEG/U13  ( .ZN(\SADR/SELSEG/n9114 ), .A(
        \SADR/SELSEG/n9094 ) );
    snl_invx2 \SADR/SELSEG/U14  ( .ZN(\SADR/SELSEG/n9107 ), .A(
        \SADR/SELSEG/n9087 ) );
    snl_invx2 \SADR/SELSEG/U21  ( .ZN(\SADR/SELSEG/n9100 ), .A(
        \SADR/SELSEG/n9078 ) );
    snl_nand04x0 \SADR/SELSEG/U54  ( .ZN(\SADR/lmtaddr[10] ), .A(
        \SADR/SELSEG/n9041 ), .B(\SADR/SELSEG/n9042 ), .C(\SADR/SELSEG/n9043 ), 
        .D(\SADR/SELSEG/n9044 ) );
    snl_nand02x1 \SADR/SELSEG/U73  ( .ZN(\SADR/SELSEG/n9082 ), .A(
        \SADR/SELSEG/n9081 ), .B(\SADR/SELSEG/n9075 ) );
    snl_aoi2222x0 \SADR/SELSEG/U113  ( .ZN(\SADR/SELSEG/n8953 ), .A(
        \pk_s3ba_h[6] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[6] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[6] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[6] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U223  ( .ZN(\SADR/SELSEG/n9047 ), .A(
        \pk_sabl_h[27] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[11] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[27] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[11] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U134  ( .ZN(\SADR/SELSEG/n9000 ), .A(
        \pk_sfba_h[17] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[17] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[17] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[17] ), .H(\SADR/SELSEG/n9102 ) );
    snl_oai2222x0 \SADR/SELSEG/U96  ( .ZN(\SADR/SELSEG/n9068 ), .A(
        \ph_segset_h[4] ), .B(\SADR/SELSEG/n9092 ), .C(\ph_segset_h[5] ), .D(
        \SADR/SELSEG/n9091 ), .E(\ph_segset_h[6] ), .F(\SADR/SELSEG/n9090 ), 
        .G(\ph_segset_h[7] ), .H(\SADR/SELSEG/n9089 ) );
    snl_aoi2222x0 \SADR/SELSEG/U198  ( .ZN(\SADR/SELSEG/n9012 ), .A(
        \pk_sefl_h[18] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[2] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[18] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[2] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U204  ( .ZN(\SADR/SELSEG/n9006 ), .A(
        \pk_s67l_h[17] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[1] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[17] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[1] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U166  ( .ZN(\SADR/SELSEG/n8932 ), .A(
        \pk_sfba_h[0] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[0] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[0] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[0] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nor02x1 \SADR/SELSEG/U68  ( .ZN(\SADR/SELSEG/n9077 ), .A(
        \SADR/SELSEG/n9073 ), .B(\pgsdprhh[28] ) );
    snl_aoi2222x0 \SADR/SELSEG/U108  ( .ZN(\SADR/SELSEG/n8958 ), .A(
        \pk_s7ba_h[7] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[7] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[7] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[7] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U141  ( .ZN(\SADR/SELSEG/n8993 ), .A(
        \pk_s3ba_h[16] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[16] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[16] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[16] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U183  ( .ZN(\SADR/SELSEG/n9027 ), .A(
        \pk_sabl_h[22] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[6] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[22] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[6] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U174  ( .ZN(\SADR/SELSEG/n9036 ), .A(
        \pk_sefl_h[24] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[8] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[24] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[8] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U191  ( .ZN(\SADR/SELSEG/n9019 ), .A(
        \pk_sabl_h[20] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[4] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[20] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[4] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nand04x0 \SADR/SELSEG/U28  ( .ZN(\SADR/segbase[2] ), .A(
        \SADR/SELSEG/n8937 ), .B(\SADR/SELSEG/n8938 ), .C(\SADR/SELSEG/n8939 ), 
        .D(\SADR/SELSEG/n8940 ) );
    snl_nand04x0 \SADR/SELSEG/U33  ( .ZN(\SADR/segbase[7] ), .A(
        \SADR/SELSEG/n8957 ), .B(\SADR/SELSEG/n8958 ), .C(\SADR/SELSEG/n8959 ), 
        .D(\SADR/SELSEG/n8960 ) );
    snl_aoi2222x0 \SADR/SELSEG/U148  ( .ZN(\SADR/SELSEG/n8986 ), .A(
        \pk_s7ba_h[14] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[14] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[14] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[14] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U153  ( .ZN(\SADR/SELSEG/n8981 ), .A(
        \pk_s3ba_h[13] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[13] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[13] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[13] ), .H(\SADR/SELSEG/n9117 ) );
    snl_nand04x0 \SADR/SELSEG/U34  ( .ZN(\SADR/segbase[8] ), .A(
        \SADR/SELSEG/n8961 ), .B(\SADR/SELSEG/n8962 ), .C(\SADR/SELSEG/n8963 ), 
        .D(\SADR/SELSEG/n8964 ) );
    snl_nand04x0 \SADR/SELSEG/U41  ( .ZN(\SADR/segbase[15] ), .A(
        \SADR/SELSEG/n8989 ), .B(\SADR/SELSEG/n8990 ), .C(\SADR/SELSEG/n8991 ), 
        .D(\SADR/SELSEG/n8992 ) );
    snl_nand04x0 \SADR/SELSEG/U46  ( .ZN(\SADR/lmtaddr[2] ), .A(
        \SADR/SELSEG/n9009 ), .B(\SADR/SELSEG/n9010 ), .C(\SADR/SELSEG/n9011 ), 
        .D(\SADR/SELSEG/n9012 ) );
    snl_invx05 \SADR/SELSEG/U61  ( .ZN(\SADR/SELSEG/n9070 ), .A(\pgsdprhh[30] 
        ) );
    snl_nor02x1 \SADR/SELSEG/U84  ( .ZN(\SADR/SELSEG/n9093 ), .A(
        \pgsdprhh[30] ), .B(\pgsdprhh[31] ) );
    snl_aoi2222x0 \SADR/SELSEG/U101  ( .ZN(\SADR/SELSEG/n8965 ), .A(
        \pk_s3ba_h[9] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[9] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[9] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[9] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U231  ( .ZN(\SADR/SELSEG/n9003 ), .A(
        \pk_sabl_h[16] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[0] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[16] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[0] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U126  ( .ZN(\SADR/SELSEG/n8940 ), .A(
        \pk_sfba_h[2] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[2] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[2] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[2] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U211  ( .ZN(\SADR/SELSEG/n9059 ), .A(
        \pk_sabl_h[30] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[14] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[30] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[14] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U216  ( .ZN(\SADR/SELSEG/n9054 ), .A(
        \pk_s67l_h[29] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[13] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[29] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[13] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nor02x1 \SADR/SELSEG/U66  ( .ZN(\SADR/SELSEG/n9075 ), .A(
        \SADR/SELSEG/n9071 ), .B(\SADR/SELSEG/n9070 ) );
    snl_aoi2222x0 \SADR/SELSEG/U106  ( .ZN(\SADR/SELSEG/n8960 ), .A(
        \pk_sfba_h[7] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[7] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[7] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[7] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U121  ( .ZN(\SADR/SELSEG/n8945 ), .A(
        \pk_s3ba_h[4] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[4] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[4] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[4] ), .H(\SADR/SELSEG/n9117 ) );
    snl_nand02x1 \SADR/SELSEG/U83  ( .ZN(\SADR/SELSEG/n9092 ), .A(
        \SADR/SELSEG/n9088 ), .B(\SADR/SELSEG/n9081 ) );
    snl_aoi2222x0 \SADR/SELSEG/U168  ( .ZN(\SADR/SELSEG/n8930 ), .A(
        \pk_s7ba_h[0] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[0] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[0] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[0] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U98  ( .ZN(\SADR/SELSEG/n8968 ), .A(
        \pk_sfba_h[9] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[9] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[9] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[9] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U154  ( .ZN(\SADR/SELSEG/n8980 ), .A(
        \pk_sfba_h[12] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[12] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[12] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[12] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nand04x0 \SADR/SELSEG/U26  ( .ZN(\SADR/segbase[0] ), .A(
        \SADR/SELSEG/n8929 ), .B(\SADR/SELSEG/n8930 ), .C(\SADR/SELSEG/n8931 ), 
        .D(\SADR/SELSEG/n8932 ) );
    snl_nand04x0 \SADR/SELSEG/U48  ( .ZN(\SADR/lmtaddr[4] ), .A(
        \SADR/SELSEG/n9017 ), .B(\SADR/SELSEG/n9018 ), .C(\SADR/SELSEG/n9019 ), 
        .D(\SADR/SELSEG/n9020 ) );
    snl_aoi2222x0 \SADR/SELSEG/U128  ( .ZN(\SADR/SELSEG/n8938 ), .A(
        \pk_s7ba_h[2] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[2] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[2] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[2] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U173  ( .ZN(\SADR/SELSEG/n9037 ), .A(
        \pk_s23l_h[25] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[9] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[25] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[9] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U184  ( .ZN(\SADR/SELSEG/n9026 ), .A(
        \pk_s67l_h[22] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[6] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[22] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[6] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U196  ( .ZN(\SADR/SELSEG/n9014 ), .A(
        \pk_s67l_h[19] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[3] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[19] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[3] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U146  ( .ZN(\SADR/SELSEG/n8988 ), .A(
        \pk_sfba_h[14] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[14] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[14] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[14] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U218  ( .ZN(\SADR/SELSEG/n9052 ), .A(
        \pk_sefl_h[28] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[12] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[28] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[12] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nand04x0 \SADR/SELSEG/U35  ( .ZN(\SADR/segbase[9] ), .A(
        \SADR/SELSEG/n8965 ), .B(\SADR/SELSEG/n8966 ), .C(\SADR/SELSEG/n8967 ), 
        .D(\SADR/SELSEG/n8968 ) );
    snl_nand04x0 \SADR/SELSEG/U53  ( .ZN(\SADR/lmtaddr[9] ), .A(
        \SADR/SELSEG/n9037 ), .B(\SADR/SELSEG/n9038 ), .C(\SADR/SELSEG/n9039 ), 
        .D(\SADR/SELSEG/n9040 ) );
    snl_aoi2222x0 \SADR/SELSEG/U91  ( .ZN(\SADR/SELSEG/n9108 ), .A(
        \SADR/SELSEG/n9109 ), .B(\ph_segset_h[23] ), .C(\SADR/SELSEG/n9110 ), 
        .D(\ph_segset_h[22] ), .E(\SADR/SELSEG/n9111 ), .F(\ph_segset_h[21] ), 
        .G(\SADR/SELSEG/n9112 ), .H(\ph_segset_h[20] ) );
    snl_aoi2222x0 \SADR/SELSEG/U161  ( .ZN(\SADR/SELSEG/n8973 ), .A(
        \pk_s3ba_h[11] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[11] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[11] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[11] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U203  ( .ZN(\SADR/SELSEG/n9007 ), .A(
        \pk_sabl_h[17] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[1] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[17] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[1] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nor02x1 \SADR/SELSEG/U74  ( .ZN(\SADR/SELSEG/n9083 ), .A(
        \SADR/SELSEG/n9071 ), .B(\pgsdprhh[30] ) );
    snl_aoi2222x0 \SADR/SELSEG/U114  ( .ZN(\SADR/SELSEG/n8952 ), .A(
        \pk_sfba_h[5] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[5] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[5] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[5] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U133  ( .ZN(\SADR/SELSEG/n8933 ), .A(
        \pk_s3ba_h[1] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[1] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[1] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[1] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U224  ( .ZN(\SADR/SELSEG/n9046 ), .A(
        \pk_s67l_h[27] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[11] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[27] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[11] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U99  ( .ZN(\SADR/SELSEG/n8967 ), .A(
        \pk_sbba_h[9] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[9] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[9] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[9] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U197  ( .ZN(\SADR/SELSEG/n9013 ), .A(
        \pk_s23l_h[19] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[3] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[19] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[3] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U155  ( .ZN(\SADR/SELSEG/n8979 ), .A(
        \pk_sbba_h[12] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[12] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[12] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[12] ), .H(\SADR/SELSEG/n9107 ) );
    snl_invx2 \SADR/SELSEG/U15  ( .ZN(\SADR/SELSEG/n9112 ), .A(
        \SADR/SELSEG/n9092 ) );
    snl_invx2 \SADR/SELSEG/U20  ( .ZN(\SADR/SELSEG/n9115 ), .A(
        \SADR/SELSEG/n9095 ) );
    snl_nand04x0 \SADR/SELSEG/U27  ( .ZN(\SADR/segbase[1] ), .A(
        \SADR/SELSEG/n8933 ), .B(\SADR/SELSEG/n8934 ), .C(\SADR/SELSEG/n8935 ), 
        .D(\SADR/SELSEG/n8936 ) );
    snl_nand04x0 \SADR/SELSEG/U40  ( .ZN(\SADR/segbase[14] ), .A(
        \SADR/SELSEG/n8985 ), .B(\SADR/SELSEG/n8986 ), .C(\SADR/SELSEG/n8987 ), 
        .D(\SADR/SELSEG/n8988 ) );
    snl_nand02x1 \SADR/SELSEG/U82  ( .ZN(\SADR/SELSEG/n9091 ), .A(
        \SADR/SELSEG/n9088 ), .B(\SADR/SELSEG/n9079 ) );
    snl_aoi2222x0 \SADR/SELSEG/U169  ( .ZN(\SADR/SELSEG/n8929 ), .A(
        \pk_s3ba_h[0] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[0] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[0] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[0] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U172  ( .ZN(\SADR/SELSEG/n9038 ), .A(
        \pk_s67l_h[25] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[9] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[25] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[9] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nand04x0 \SADR/SELSEG/U52  ( .ZN(\SADR/lmtaddr[8] ), .A(
        \SADR/SELSEG/n9033 ), .B(\SADR/SELSEG/n9034 ), .C(\SADR/SELSEG/n9035 ), 
        .D(\SADR/SELSEG/n9036 ) );
    snl_nand02x1 \SADR/SELSEG/U67  ( .ZN(\SADR/SELSEG/n9076 ), .A(
        \SADR/SELSEG/n9075 ), .B(\SADR/SELSEG/n9074 ) );
    snl_aoi2222x0 \SADR/SELSEG/U107  ( .ZN(\SADR/SELSEG/n8959 ), .A(
        \pk_sbba_h[7] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[7] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[7] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[7] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U120  ( .ZN(\SADR/SELSEG/n8946 ), .A(
        \pk_s7ba_h[4] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[4] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[4] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[4] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U210  ( .ZN(\SADR/SELSEG/n9060 ), .A(
        \pk_sefl_h[30] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[14] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[30] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[14] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nand02x1 \SADR/SELSEG/U75  ( .ZN(\SADR/SELSEG/n9084 ), .A(
        \SADR/SELSEG/n9083 ), .B(\SADR/SELSEG/n9074 ) );
    snl_aoi2222x0 \SADR/SELSEG/U115  ( .ZN(\SADR/SELSEG/n8951 ), .A(
        \pk_sbba_h[5] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[5] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[5] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[5] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U132  ( .ZN(\SADR/SELSEG/n8934 ), .A(
        \pk_s7ba_h[1] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[1] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[1] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[1] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U202  ( .ZN(\SADR/SELSEG/n9008 ), .A(
        \pk_sefl_h[17] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[1] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[17] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[1] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U90  ( .ZN(\SADR/SELSEG/n9103 ), .A(
        \SADR/SELSEG/n9104 ), .B(\ph_segset_h[27] ), .C(\SADR/SELSEG/n9105 ), 
        .D(\ph_segset_h[26] ), .E(\SADR/SELSEG/n9106 ), .F(\ph_segset_h[25] ), 
        .G(\SADR/SELSEG/n9107 ), .H(\ph_segset_h[24] ) );
    snl_aoi2222x0 \SADR/SELSEG/U225  ( .ZN(\SADR/SELSEG/n9045 ), .A(
        \pk_s23l_h[27] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[11] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[27] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[11] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U147  ( .ZN(\SADR/SELSEG/n8987 ), .A(
        \pk_sbba_h[14] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[14] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[14] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[14] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nand04x0 \SADR/SELSEG/U49  ( .ZN(\SADR/lmtaddr[5] ), .A(
        \SADR/SELSEG/n9021 ), .B(\SADR/SELSEG/n9022 ), .C(\SADR/SELSEG/n9023 ), 
        .D(\SADR/SELSEG/n9024 ) );
    snl_aoi2222x0 \SADR/SELSEG/U129  ( .ZN(\SADR/SELSEG/n8937 ), .A(
        \pk_s3ba_h[2] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[2] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[2] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[2] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U160  ( .ZN(\SADR/SELSEG/n8974 ), .A(
        \pk_s7ba_h[11] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[11] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[11] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[11] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U185  ( .ZN(\SADR/SELSEG/n9025 ), .A(
        \pk_s23l_h[22] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[6] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[22] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[6] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U219  ( .ZN(\SADR/SELSEG/n9051 ), .A(
        \pk_sabl_h[28] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[12] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[28] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[12] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nand02x1 \SADR/SELSEG/U69  ( .ZN(\SADR/SELSEG/n9078 ), .A(
        \SADR/SELSEG/n9077 ), .B(\SADR/SELSEG/n9075 ) );
    snl_aoi2222x0 \SADR/SELSEG/U109  ( .ZN(\SADR/SELSEG/n8957 ), .A(
        \pk_s3ba_h[7] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[7] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[7] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[7] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U182  ( .ZN(\SADR/SELSEG/n9028 ), .A(
        \pk_sefl_h[22] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[6] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[22] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[6] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U167  ( .ZN(\SADR/SELSEG/n8931 ), .A(
        \pk_sbba_h[0] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[0] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[0] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[0] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nand04x0 \SADR/SELSEG/U29  ( .ZN(\SADR/segbase[3] ), .A(
        \SADR/SELSEG/n8941 ), .B(\SADR/SELSEG/n8942 ), .C(\SADR/SELSEG/n8943 ), 
        .D(\SADR/SELSEG/n8944 ) );
    snl_nand04x0 \SADR/SELSEG/U47  ( .ZN(\SADR/lmtaddr[3] ), .A(
        \SADR/SELSEG/n9013 ), .B(\SADR/SELSEG/n9014 ), .C(\SADR/SELSEG/n9015 ), 
        .D(\SADR/SELSEG/n9016 ) );
    snl_nand04x0 \SADR/SELSEG/U55  ( .ZN(\SADR/lmtaddr[11] ), .A(
        \SADR/SELSEG/n9045 ), .B(\SADR/SELSEG/n9046 ), .C(\SADR/SELSEG/n9047 ), 
        .D(\SADR/SELSEG/n9048 ) );
    snl_nor02x1 \SADR/SELSEG/U72  ( .ZN(\SADR/SELSEG/n9081 ), .A(
        \pgsdprhh[28] ), .B(\pgsdprhh[29] ) );
    snl_oai2222x0 \SADR/SELSEG/U97  ( .ZN(\SADR/SELSEG/n9069 ), .A(
        \ph_segset_h[0] ), .B(\SADR/SELSEG/n9097 ), .C(\ph_segset_h[1] ), .D(
        \SADR/SELSEG/n9096 ), .E(\ph_segset_h[2] ), .F(\SADR/SELSEG/n9095 ), 
        .G(\ph_segset_h[3] ), .H(\SADR/SELSEG/n9094 ) );
    snl_aoi2222x0 \SADR/SELSEG/U140  ( .ZN(\SADR/SELSEG/n8994 ), .A(
        \pk_s7ba_h[16] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[16] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[16] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[16] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U222  ( .ZN(\SADR/SELSEG/n9048 ), .A(
        \pk_sefl_h[27] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[11] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[27] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[11] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U112  ( .ZN(\SADR/SELSEG/n8954 ), .A(
        \pk_s7ba_h[6] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[6] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[6] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[6] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U135  ( .ZN(\SADR/SELSEG/n8999 ), .A(
        \pk_sbba_h[17] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[17] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[17] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[17] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U205  ( .ZN(\SADR/SELSEG/n9005 ), .A(
        \pk_s23l_h[17] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[1] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[17] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[1] ), .H(\SADR/SELSEG/n9117 ) );
    snl_or05x1 \SADR/SELSEG/U60  ( .Z(\SADR/seglmterr ), .A(
        \SADR/SELSEG/n9065 ), .B(\SADR/SELSEG/n9066 ), .C(\SADR/SELSEG/n9067 ), 
        .D(\SADR/SELSEG/n9068 ), .E(\SADR/SELSEG/n9069 ) );
    snl_aoi2222x0 \SADR/SELSEG/U199  ( .ZN(\SADR/SELSEG/n9011 ), .A(
        \pk_sabl_h[18] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[2] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[18] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[2] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U230  ( .ZN(\SADR/SELSEG/n9004 ), .A(
        \pk_sefl_h[16] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[0] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[16] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[0] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U100  ( .ZN(\SADR/SELSEG/n8966 ), .A(
        \pk_s7ba_h[9] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[9] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[9] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[9] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U127  ( .ZN(\SADR/SELSEG/n8939 ), .A(
        \pk_sbba_h[2] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[2] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[2] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[2] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U217  ( .ZN(\SADR/SELSEG/n9053 ), .A(
        \pk_s23l_h[29] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[13] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[29] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[13] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U149  ( .ZN(\SADR/SELSEG/n8985 ), .A(
        \pk_s3ba_h[14] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[14] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[14] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[14] ), .H(\SADR/SELSEG/n9117 ) );
    snl_nand02x1 \SADR/SELSEG/U85  ( .ZN(\SADR/SELSEG/n9094 ), .A(
        \SADR/SELSEG/n9093 ), .B(\SADR/SELSEG/n9074 ) );
    snl_aoi2222x0 \SADR/SELSEG/U175  ( .ZN(\SADR/SELSEG/n9035 ), .A(
        \pk_sabl_h[24] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[8] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[24] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[8] ), .H(\SADR/SELSEG/n9107 ) );
    snl_invx2 \SADR/SELSEG/U17  ( .ZN(\SADR/SELSEG/n9117 ), .A(
        \SADR/SELSEG/n9097 ) );
    snl_invx2 \SADR/SELSEG/U22  ( .ZN(\SADR/SELSEG/n9111 ), .A(
        \SADR/SELSEG/n9091 ) );
    snl_nand04x0 \SADR/SELSEG/U32  ( .ZN(\SADR/segbase[6] ), .A(
        \SADR/SELSEG/n8953 ), .B(\SADR/SELSEG/n8954 ), .C(\SADR/SELSEG/n8955 ), 
        .D(\SADR/SELSEG/n8956 ) );
    snl_nand04x0 \SADR/SELSEG/U39  ( .ZN(\SADR/segbase[13] ), .A(
        \SADR/SELSEG/n8981 ), .B(\SADR/SELSEG/n8982 ), .C(\SADR/SELSEG/n8983 ), 
        .D(\SADR/SELSEG/n8984 ) );
    snl_nand04x0 \SADR/SELSEG/U57  ( .ZN(\SADR/lmtaddr[13] ), .A(
        \SADR/SELSEG/n9053 ), .B(\SADR/SELSEG/n9054 ), .C(\SADR/SELSEG/n9055 ), 
        .D(\SADR/SELSEG/n9056 ) );
    snl_aoi2222x0 \SADR/SELSEG/U137  ( .ZN(\SADR/SELSEG/n8997 ), .A(
        \pk_s3ba_h[17] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[17] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[17] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[17] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U152  ( .ZN(\SADR/SELSEG/n8982 ), .A(
        \pk_s7ba_h[13] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[13] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[13] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[13] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U190  ( .ZN(\SADR/SELSEG/n9020 ), .A(
        \pk_sefl_h[20] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[4] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[20] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[4] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nor02x1 \SADR/SELSEG/U70  ( .ZN(\SADR/SELSEG/n9079 ), .A(
        \SADR/SELSEG/n9072 ), .B(\pgsdprhh[29] ) );
    snl_aoi2222x0 \SADR/SELSEG/U207  ( .ZN(\SADR/SELSEG/n9063 ), .A(
        \pk_sabl_h[31] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[15] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[31] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[15] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U110  ( .ZN(\SADR/SELSEG/n8956 ), .A(
        \pk_sfba_h[6] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[6] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[6] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[6] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U220  ( .ZN(\SADR/SELSEG/n9050 ), .A(
        \pk_s67l_h[28] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[12] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[28] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[12] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U159  ( .ZN(\SADR/SELSEG/n8975 ), .A(
        \pk_sbba_h[11] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[11] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[11] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[11] ), .H(\SADR/SELSEG/n9107 ) );
    snl_oai2222x0 \SADR/SELSEG/U95  ( .ZN(\SADR/SELSEG/n9067 ), .A(
        \ph_segset_h[8] ), .B(\SADR/SELSEG/n9087 ), .C(\ph_segset_h[9] ), .D(
        \SADR/SELSEG/n9086 ), .E(\ph_segset_h[10] ), .F(\SADR/SELSEG/n9085 ), 
        .G(\ph_segset_h[11] ), .H(\SADR/SELSEG/n9084 ) );
    snl_nand04x0 \SADR/SELSEG/U30  ( .ZN(\SADR/segbase[4] ), .A(
        \SADR/SELSEG/n8945 ), .B(\SADR/SELSEG/n8946 ), .C(\SADR/SELSEG/n8947 ), 
        .D(\SADR/SELSEG/n8948 ) );
    snl_nor02x1 \SADR/SELSEG/U79  ( .ZN(\SADR/SELSEG/n9088 ), .A(
        \SADR/SELSEG/n9070 ), .B(\pgsdprhh[31] ) );
    snl_aoi2222x0 \SADR/SELSEG/U119  ( .ZN(\SADR/SELSEG/n8947 ), .A(
        \pk_sbba_h[4] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[4] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[4] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[4] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U142  ( .ZN(\SADR/SELSEG/n8992 ), .A(
        \pk_sfba_h[15] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[15] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[15] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[15] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U165  ( .ZN(\SADR/SELSEG/n8969 ), .A(
        \pk_s3ba_h[10] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[10] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[10] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[10] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U180  ( .ZN(\SADR/SELSEG/n9030 ), .A(
        \pk_s67l_h[23] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[7] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[23] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[7] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U192  ( .ZN(\SADR/SELSEG/n9018 ), .A(
        \pk_s67l_h[20] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[4] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[20] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[4] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U229  ( .ZN(\SADR/SELSEG/n9041 ), .A(
        \pk_s23l_h[26] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[10] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[26] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[10] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U150  ( .ZN(\SADR/SELSEG/n8984 ), .A(
        \pk_sfba_h[13] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[13] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[13] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[13] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U177  ( .ZN(\SADR/SELSEG/n9033 ), .A(
        \pk_s23l_h[24] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[8] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[24] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[8] ), .H(\SADR/SELSEG/n9117 ) );
    snl_nand04x0 \SADR/SELSEG/U42  ( .ZN(\SADR/segbase[16] ), .A(
        \SADR/SELSEG/n8993 ), .B(\SADR/SELSEG/n8994 ), .C(\SADR/SELSEG/n8995 ), 
        .D(\SADR/SELSEG/n8996 ) );
    snl_nand04x0 \SADR/SELSEG/U45  ( .ZN(\SADR/lmtaddr[1] ), .A(
        \SADR/SELSEG/n9005 ), .B(\SADR/SELSEG/n9006 ), .C(\SADR/SELSEG/n9007 ), 
        .D(\SADR/SELSEG/n9008 ) );
    snl_nand02x1 \SADR/SELSEG/U87  ( .ZN(\SADR/SELSEG/n9096 ), .A(
        \SADR/SELSEG/n9093 ), .B(\SADR/SELSEG/n9079 ) );
    snl_aoi2222x0 \SADR/SELSEG/U125  ( .ZN(\SADR/SELSEG/n8941 ), .A(
        \pk_s3ba_h[3] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[3] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[3] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[3] ), .H(\SADR/SELSEG/n9117 ) );
    snl_invx05 \SADR/SELSEG/U62  ( .ZN(\SADR/SELSEG/n9071 ), .A(\pgsdprhh[31] 
        ) );
    snl_aoi2222x0 \SADR/SELSEG/U215  ( .ZN(\SADR/SELSEG/n9055 ), .A(
        \pk_sabl_h[29] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[13] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[29] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[13] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nor02x1 \SADR/SELSEG/U65  ( .ZN(\SADR/SELSEG/n9074 ), .A(
        \SADR/SELSEG/n9073 ), .B(\SADR/SELSEG/n9072 ) );
    snl_aoi2222x0 \SADR/SELSEG/U102  ( .ZN(\SADR/SELSEG/n8964 ), .A(
        \pk_sfba_h[8] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[8] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[8] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[8] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U232  ( .ZN(\SADR/SELSEG/n9002 ), .A(
        \pk_s67l_h[16] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[0] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[16] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[0] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U105  ( .ZN(\SADR/SELSEG/n8961 ), .A(
        \pk_s3ba_h[8] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[8] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[8] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[8] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U189  ( .ZN(\SADR/SELSEG/n9021 ), .A(
        \pk_s23l_h[21] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[5] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[21] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[5] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U212  ( .ZN(\SADR/SELSEG/n9058 ), .A(
        \pk_s67l_h[30] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[14] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[30] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[14] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nand02x1 \SADR/SELSEG/U80  ( .ZN(\SADR/SELSEG/n9089 ), .A(
        \SADR/SELSEG/n9088 ), .B(\SADR/SELSEG/n9074 ) );
    snl_aoi2222x0 \SADR/SELSEG/U122  ( .ZN(\SADR/SELSEG/n8944 ), .A(
        \pk_sfba_h[3] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[3] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[3] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[3] ), .H(\SADR/SELSEG/n9102 ) );
    snl_invx1 \SADR/SELSEG/U11  ( .ZN(\SADR/SELSEG/n9109 ), .A(
        \SADR/SELSEG/n9089 ) );
    snl_invx2 \SADR/SELSEG/U19  ( .ZN(\SADR/SELSEG/n9105 ), .A(
        \SADR/SELSEG/n9085 ) );
    snl_invx2 \SADR/SELSEG/U25  ( .ZN(\SADR/SELSEG/n9101 ), .A(
        \SADR/SELSEG/n9080 ) );
    snl_nand04x0 \SADR/SELSEG/U37  ( .ZN(\SADR/segbase[11] ), .A(
        \SADR/SELSEG/n8973 ), .B(\SADR/SELSEG/n8974 ), .C(\SADR/SELSEG/n8975 ), 
        .D(\SADR/SELSEG/n8976 ) );
    snl_aoi2222x0 \SADR/SELSEG/U157  ( .ZN(\SADR/SELSEG/n8977 ), .A(
        \pk_s3ba_h[12] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[12] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[12] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[12] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U170  ( .ZN(\SADR/SELSEG/n9040 ), .A(
        \pk_sefl_h[25] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[9] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[25] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[9] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nand04x0 \SADR/SELSEG/U59  ( .ZN(\SADR/lmtaddr[15] ), .A(
        \SADR/SELSEG/n9061 ), .B(\SADR/SELSEG/n9062 ), .C(\SADR/SELSEG/n9063 ), 
        .D(\SADR/SELSEG/n9064 ) );
    snl_aoi2222x0 \SADR/SELSEG/U139  ( .ZN(\SADR/SELSEG/n8995 ), .A(
        \pk_sbba_h[16] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[16] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[16] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[16] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U195  ( .ZN(\SADR/SELSEG/n9015 ), .A(
        \pk_sabl_h[19] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[3] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[19] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[3] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U89  ( .ZN(\SADR/SELSEG/n9098 ), .A(
        \SADR/SELSEG/n9099 ), .B(\ph_segset_h[31] ), .C(\SADR/SELSEG/n9100 ), 
        .D(\ph_segset_h[30] ), .E(\SADR/SELSEG/n9101 ), .F(\ph_segset_h[29] ), 
        .G(\SADR/SELSEG/n9102 ), .H(\ph_segset_h[28] ) );
    snl_aoi2222x0 \SADR/SELSEG/U187  ( .ZN(\SADR/SELSEG/n9023 ), .A(
        \pk_sabl_h[21] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[5] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[21] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[5] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U209  ( .ZN(\SADR/SELSEG/n9061 ), .A(
        \pk_s23l_h[31] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[15] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[31] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[15] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U145  ( .ZN(\SADR/SELSEG/n8989 ), .A(
        \pk_s3ba_h[15] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[15] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[15] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s0ba_h[15] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U162  ( .ZN(\SADR/SELSEG/n8972 ), .A(
        \pk_sfba_h[10] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[10] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[10] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[10] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U179  ( .ZN(\SADR/SELSEG/n9031 ), .A(
        \pk_sabl_h[23] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[7] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[23] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[7] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nand04x0 \SADR/SELSEG/U50  ( .ZN(\SADR/lmtaddr[6] ), .A(
        \SADR/SELSEG/n9025 ), .B(\SADR/SELSEG/n9026 ), .C(\SADR/SELSEG/n9027 ), 
        .D(\SADR/SELSEG/n9028 ) );
    snl_nand02x1 \SADR/SELSEG/U77  ( .ZN(\SADR/SELSEG/n9086 ), .A(
        \SADR/SELSEG/n9083 ), .B(\SADR/SELSEG/n9079 ) );
    snl_aoi2222x0 \SADR/SELSEG/U92  ( .ZN(\SADR/SELSEG/n9113 ), .A(
        \SADR/SELSEG/n9114 ), .B(\ph_segset_h[19] ), .C(\SADR/SELSEG/n9115 ), 
        .D(\ph_segset_h[18] ), .E(\SADR/SELSEG/n9116 ), .F(\ph_segset_h[17] ), 
        .G(\SADR/SELSEG/n9117 ), .H(\ph_segset_h[16] ) );
    snl_aoi2222x0 \SADR/SELSEG/U117  ( .ZN(\SADR/SELSEG/n8949 ), .A(
        \pk_s3ba_h[5] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s2ba_h[5] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s1ba_h[5] ), .F(\SADR/SELSEG/n9116 ), .G(
        \pk_s0ba_h[5] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U227  ( .ZN(\SADR/SELSEG/n9043 ), .A(
        \pk_sabl_h[26] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[10] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[26] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[10] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U200  ( .ZN(\SADR/SELSEG/n9010 ), .A(
        \pk_s67l_h[18] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[2] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[18] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[2] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nand04x0 \SADR/SELSEG/U58  ( .ZN(\SADR/lmtaddr[14] ), .A(
        \SADR/SELSEG/n9057 ), .B(\SADR/SELSEG/n9058 ), .C(\SADR/SELSEG/n9059 ), 
        .D(\SADR/SELSEG/n9060 ) );
    snl_aoi2222x0 \SADR/SELSEG/U130  ( .ZN(\SADR/SELSEG/n8936 ), .A(
        \pk_sfba_h[1] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[1] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[1] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[1] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U138  ( .ZN(\SADR/SELSEG/n8996 ), .A(
        \pk_sfba_h[16] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[16] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[16] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[16] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U194  ( .ZN(\SADR/SELSEG/n9016 ), .A(
        \pk_sefl_h[19] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[3] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[19] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[3] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U208  ( .ZN(\SADR/SELSEG/n9062 ), .A(
        \pk_s67l_h[31] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[15] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[31] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[15] ), .H(\SADR/SELSEG/n9112 ) );
    snl_invx2 \SADR/SELSEG/U16  ( .ZN(\SADR/SELSEG/n9102 ), .A(
        \SADR/SELSEG/n9082 ) );
    snl_invx2 \SADR/SELSEG/U18  ( .ZN(\SADR/SELSEG/n9110 ), .A(
        \SADR/SELSEG/n9090 ) );
    snl_nand04x0 \SADR/SELSEG/U36  ( .ZN(\SADR/segbase[10] ), .A(
        \SADR/SELSEG/n8969 ), .B(\SADR/SELSEG/n8970 ), .C(\SADR/SELSEG/n8971 ), 
        .D(\SADR/SELSEG/n8972 ) );
    snl_aoi2222x0 \SADR/SELSEG/U156  ( .ZN(\SADR/SELSEG/n8978 ), .A(
        \pk_s7ba_h[12] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[12] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[12] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[12] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U171  ( .ZN(\SADR/SELSEG/n9039 ), .A(
        \pk_sabl_h[25] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_sabl_h[9] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s89l_h[25] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s89l_h[9] ), .H(\SADR/SELSEG/n9107 ) );
    snl_nand04x0 \SADR/SELSEG/U43  ( .ZN(\SADR/segbase[17] ), .A(
        \SADR/SELSEG/n8997 ), .B(\SADR/SELSEG/n8998 ), .C(\SADR/SELSEG/n8999 ), 
        .D(\SADR/SELSEG/n9000 ) );
    snl_invx05 \SADR/SELSEG/U64  ( .ZN(\SADR/SELSEG/n9073 ), .A(\pgsdprhh[29] 
        ) );
    snl_nand02x1 \SADR/SELSEG/U81  ( .ZN(\SADR/SELSEG/n9090 ), .A(
        \SADR/SELSEG/n9088 ), .B(\SADR/SELSEG/n9077 ) );
    snl_aoi2222x0 \SADR/SELSEG/U104  ( .ZN(\SADR/SELSEG/n8962 ), .A(
        \pk_s7ba_h[8] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[8] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[8] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[8] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nand04x0 \SADR/SELSEG/U234  ( .ZN(\SADR/SELSEG/n9118 ), .A(
        \SADR/SELSEG/n9113 ), .B(\SADR/SELSEG/n9108 ), .C(\SADR/SELSEG/n9103 ), 
        .D(\SADR/SELSEG/n9098 ) );
    snl_nand04x0 \SADR/SELSEG/U51  ( .ZN(\SADR/lmtaddr[7] ), .A(
        \SADR/SELSEG/n9029 ), .B(\SADR/SELSEG/n9030 ), .C(\SADR/SELSEG/n9031 ), 
        .D(\SADR/SELSEG/n9032 ) );
    snl_nand02x1 \SADR/SELSEG/U76  ( .ZN(\SADR/SELSEG/n9085 ), .A(
        \SADR/SELSEG/n9083 ), .B(\SADR/SELSEG/n9077 ) );
    snl_aoi2222x0 \SADR/SELSEG/U116  ( .ZN(\SADR/SELSEG/n8950 ), .A(
        \pk_s7ba_h[5] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[5] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[5] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[5] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U123  ( .ZN(\SADR/SELSEG/n8943 ), .A(
        \pk_sbba_h[3] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[3] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[3] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[3] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U213  ( .ZN(\SADR/SELSEG/n9057 ), .A(
        \pk_s23l_h[30] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[14] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[30] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[14] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U226  ( .ZN(\SADR/SELSEG/n9044 ), .A(
        \pk_sefl_h[26] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[10] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[26] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[10] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U131  ( .ZN(\SADR/SELSEG/n8935 ), .A(
        \pk_sbba_h[1] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[1] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[1] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[1] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U201  ( .ZN(\SADR/SELSEG/n9009 ), .A(
        \pk_s23l_h[18] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[2] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[18] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[2] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U178  ( .ZN(\SADR/SELSEG/n9032 ), .A(
        \pk_sefl_h[23] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[7] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[23] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[7] ), .H(\SADR/SELSEG/n9102 ) );
    snl_invx2 \SADR/SELSEG/U23  ( .ZN(\SADR/SELSEG/n9106 ), .A(
        \SADR/SELSEG/n9086 ) );
    snl_invx2 \SADR/SELSEG/U24  ( .ZN(\SADR/SELSEG/n9116 ), .A(
        \SADR/SELSEG/n9096 ) );
    snl_nand02x1 \SADR/SELSEG/U88  ( .ZN(\SADR/SELSEG/n9097 ), .A(
        \SADR/SELSEG/n9093 ), .B(\SADR/SELSEG/n9081 ) );
    snl_ao2b2b2x0 \SADR/SELSEG/U93  ( .Z(\SADR/SELSEG/n9065 ), .A(
        \ph_segset_h[15] ), .B(\SADR/SELSEG/n9076 ), .C(\ph_segset_h[14] ), 
        .D(\SADR/SELSEG/n9078 ), .E(ph_atchkenh), .F(\SADR/SELSEG/n9118 ) );
    snl_aoi2222x0 \SADR/SELSEG/U144  ( .ZN(\SADR/SELSEG/n8990 ), .A(
        \pk_s7ba_h[15] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[15] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[15] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[15] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U163  ( .ZN(\SADR/SELSEG/n8971 ), .A(
        \pk_sbba_h[10] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[10] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[10] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[10] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U181  ( .ZN(\SADR/SELSEG/n9029 ), .A(
        \pk_s23l_h[23] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[7] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[23] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[7] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U186  ( .ZN(\SADR/SELSEG/n9024 ), .A(
        \pk_sefl_h[21] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[5] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[21] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[5] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nand04x0 \SADR/SELSEG/U31  ( .ZN(\SADR/segbase[5] ), .A(
        \SADR/SELSEG/n8949 ), .B(\SADR/SELSEG/n8950 ), .C(\SADR/SELSEG/n8951 ), 
        .D(\SADR/SELSEG/n8952 ) );
    snl_nand04x0 \SADR/SELSEG/U38  ( .ZN(\SADR/segbase[12] ), .A(
        \SADR/SELSEG/n8977 ), .B(\SADR/SELSEG/n8978 ), .C(\SADR/SELSEG/n8979 ), 
        .D(\SADR/SELSEG/n8980 ) );
    snl_aoi2222x0 \SADR/SELSEG/U143  ( .ZN(\SADR/SELSEG/n8991 ), .A(
        \pk_sbba_h[15] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[15] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[15] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[15] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U158  ( .ZN(\SADR/SELSEG/n8976 ), .A(
        \pk_sfba_h[11] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[11] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[11] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scba_h[11] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U164  ( .ZN(\SADR/SELSEG/n8970 ), .A(
        \pk_s7ba_h[10] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[10] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[10] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[10] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nand04x0 \SADR/SELSEG/U44  ( .ZN(\SADR/lmtaddr[0] ), .A(
        \SADR/SELSEG/n9001 ), .B(\SADR/SELSEG/n9002 ), .C(\SADR/SELSEG/n9003 ), 
        .D(\SADR/SELSEG/n9004 ) );
    snl_nand04x0 \SADR/SELSEG/U56  ( .ZN(\SADR/lmtaddr[12] ), .A(
        \SADR/SELSEG/n9049 ), .B(\SADR/SELSEG/n9050 ), .C(\SADR/SELSEG/n9051 ), 
        .D(\SADR/SELSEG/n9052 ) );
    snl_oai022x1 \SADR/SELSEG/U94  ( .ZN(\SADR/SELSEG/n9066 ), .A(
        \ph_segset_h[12] ), .B(\SADR/SELSEG/n9082 ), .C(\ph_segset_h[13] ), 
        .D(\SADR/SELSEG/n9080 ) );
    snl_aoi2222x0 \SADR/SELSEG/U136  ( .ZN(\SADR/SELSEG/n8998 ), .A(
        \pk_s7ba_h[17] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[17] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[17] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s4ba_h[17] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U206  ( .ZN(\SADR/SELSEG/n9064 ), .A(
        \pk_sefl_h[31] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[15] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[31] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[15] ), .H(\SADR/SELSEG/n9102 ) );
    snl_nand02x1 \SADR/SELSEG/U71  ( .ZN(\SADR/SELSEG/n9080 ), .A(
        \SADR/SELSEG/n9079 ), .B(\SADR/SELSEG/n9075 ) );
    snl_aoi2222x0 \SADR/SELSEG/U221  ( .ZN(\SADR/SELSEG/n9049 ), .A(
        \pk_s23l_h[28] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[12] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[28] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[12] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U111  ( .ZN(\SADR/SELSEG/n8955 ), .A(
        \pk_sbba_h[6] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[6] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[6] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[6] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U124  ( .ZN(\SADR/SELSEG/n8942 ), .A(
        \pk_s7ba_h[3] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s6ba_h[3] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s5ba_h[3] ), .F(\SADR/SELSEG/n9111 ), .G(
        \pk_s4ba_h[3] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U214  ( .ZN(\SADR/SELSEG/n9056 ), .A(
        \pk_sefl_h[29] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_sefl_h[13] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_scdl_h[29] ), .F(\SADR/SELSEG/n9101 ), 
        .G(\pk_scdl_h[13] ), .H(\SADR/SELSEG/n9102 ) );
    snl_invx05 \SADR/SELSEG/U63  ( .ZN(\SADR/SELSEG/n9072 ), .A(\pgsdprhh[28] 
        ) );
    snl_aoi2222x0 \SADR/SELSEG/U233  ( .ZN(\SADR/SELSEG/n9001 ), .A(
        \pk_s23l_h[16] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[0] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[16] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[0] ), .H(\SADR/SELSEG/n9117 ) );
    snl_nand02x1 \SADR/SELSEG/U86  ( .ZN(\SADR/SELSEG/n9095 ), .A(
        \SADR/SELSEG/n9093 ), .B(\SADR/SELSEG/n9077 ) );
    snl_aoi2222x0 \SADR/SELSEG/U103  ( .ZN(\SADR/SELSEG/n8963 ), .A(
        \pk_sbba_h[8] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[8] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[8] ), .F(\SADR/SELSEG/n9106 ), .G(
        \pk_s8ba_h[8] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U188  ( .ZN(\SADR/SELSEG/n9022 ), .A(
        \pk_s67l_h[21] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[5] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[21] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[5] ), .H(\SADR/SELSEG/n9112 ) );
    snl_aoi2222x0 \SADR/SELSEG/U151  ( .ZN(\SADR/SELSEG/n8983 ), .A(
        \pk_sbba_h[13] ), .B(\SADR/SELSEG/n9104 ), .C(\pk_saba_h[13] ), .D(
        \SADR/SELSEG/n9105 ), .E(\pk_s9ba_h[13] ), .F(\SADR/SELSEG/n9106 ), 
        .G(\pk_s8ba_h[13] ), .H(\SADR/SELSEG/n9107 ) );
    snl_aoi2222x0 \SADR/SELSEG/U176  ( .ZN(\SADR/SELSEG/n9034 ), .A(
        \pk_s67l_h[24] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[8] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[24] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[8] ), .H(\SADR/SELSEG/n9112 ) );
    snl_nand02x1 \SADR/SELSEG/U78  ( .ZN(\SADR/SELSEG/n9087 ), .A(
        \SADR/SELSEG/n9083 ), .B(\SADR/SELSEG/n9081 ) );
    snl_aoi2222x0 \SADR/SELSEG/U118  ( .ZN(\SADR/SELSEG/n8948 ), .A(
        \pk_sfba_h[4] ), .B(\SADR/SELSEG/n9099 ), .C(\pk_seba_h[4] ), .D(
        \SADR/SELSEG/n9100 ), .E(\pk_sdba_h[4] ), .F(\SADR/SELSEG/n9101 ), .G(
        \pk_scba_h[4] ), .H(\SADR/SELSEG/n9102 ) );
    snl_aoi2222x0 \SADR/SELSEG/U193  ( .ZN(\SADR/SELSEG/n9017 ), .A(
        \pk_s23l_h[20] ), .B(\SADR/SELSEG/n9114 ), .C(\pk_s23l_h[4] ), .D(
        \SADR/SELSEG/n9115 ), .E(\pk_s01l_h[20] ), .F(\SADR/SELSEG/n9116 ), 
        .G(\pk_s01l_h[4] ), .H(\SADR/SELSEG/n9117 ) );
    snl_aoi2222x0 \SADR/SELSEG/U228  ( .ZN(\SADR/SELSEG/n9042 ), .A(
        \pk_s67l_h[26] ), .B(\SADR/SELSEG/n9109 ), .C(\pk_s67l_h[10] ), .D(
        \SADR/SELSEG/n9110 ), .E(\pk_s45l_h[26] ), .F(\SADR/SELSEG/n9111 ), 
        .G(\pk_s45l_h[10] ), .H(\SADR/SELSEG/n9112 ) );
    snl_ao012x1 \REG_2/ph4dec2_1/U6  ( .Z(\REG_2/ncnt3[1] ), .A(
        \REG_2/RETCNT[6] ), .B(\REG_2/RETCNT[7] ), .C(ph_errtendh) );
    snl_invx05 \REG_2/ph4dec2_1/U7  ( .ZN(\REG_2/ncnt3[0] ), .A(
        \REG_2/RETCNT[6] ) );
    snl_nor02x1 \REG_2/ph4dec2_1/U8  ( .ZN(ph_errtendh), .A(\REG_2/RETCNT[7] ), 
        .B(\REG_2/RETCNT[6] ) );
    snl_and02x1 \LBUS/ldoecnt_4/U8  ( .Z(ph_ldaoutenh4), .A(ph_lbwrh), .B(
        \LBUS/temp[3] ) );
    snl_invx05 \REGF/pbmemcnt1/add_53/U5  ( .ZN(
        \REGF/pbmemcnt1/upcnt_data283[0] ), .A(\REGF/pbmemcnt1/upcnt_data[0] )
         );
    snl_xor2x0 \REGF/pbmemcnt1/add_53/U6  ( .Z(
        \REGF/pbmemcnt1/upcnt_data283[11] ), .A(
        \REGF/pbmemcnt1/upcnt_data[11] ), .B(\REGF/pbmemcnt1/add_53/carry[11] 
        ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_10  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[10] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[11] ), .A(\REGF/pbmemcnt1/upcnt_data[10] 
        ), .B(\REGF/pbmemcnt1/add_53/carry[10] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_3  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[3] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[4] ), .A(\REGF/pbmemcnt1/upcnt_data[3] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[3] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_4  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[4] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[5] ), .A(\REGF/pbmemcnt1/upcnt_data[4] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[4] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_2  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[2] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[3] ), .A(\REGF/pbmemcnt1/upcnt_data[2] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[2] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_5  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[5] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[6] ), .A(\REGF/pbmemcnt1/upcnt_data[5] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[5] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_7  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[7] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[8] ), .A(\REGF/pbmemcnt1/upcnt_data[7] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[7] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_1  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[1] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[2] ), .A(\REGF/pbmemcnt1/upcnt_data[1] ), 
        .B(\REGF/pbmemcnt1/upcnt_data[0] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_9  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[9] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[10] ), .A(\REGF/pbmemcnt1/upcnt_data[9] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[9] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_6  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[6] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[7] ), .A(\REGF/pbmemcnt1/upcnt_data[6] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[6] ) );
    snl_add05x1 \REGF/pbmemcnt1/add_53/U1_1_8  ( .S(
        \REGF/pbmemcnt1/upcnt_data283[8] ), .CO(
        \REGF/pbmemcnt1/add_53/carry[9] ), .A(\REGF/pbmemcnt1/upcnt_data[8] ), 
        .B(\REGF/pbmemcnt1/add_53/carry[8] ) );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U6  ( .ZN(
        \REGF/pbmemcnt1/down_data274[7] ), .A(\REGF/pbmemcnt1/down_data[7] ), 
        .B(\REGF/pbmemcnt1/sub_48/carry[7] ) );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U14  ( .ZN(
        \REGF/pbmemcnt1/down_data274[3] ), .A(\REGF/pbmemcnt1/sub_48/carry[3] 
        ), .B(\REGF/pbmemcnt1/down_data[3] ) );
    snl_or02x1 \REGF/pbmemcnt1/sub_48/U7  ( .Z(
        \REGF/pbmemcnt1/sub_48/carry[7] ), .A(\REGF/pbmemcnt1/down_data[6] ), 
        .B(\REGF/pbmemcnt1/sub_48/carry[6] ) );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U8  ( .ZN(
        \REGF/pbmemcnt1/down_data274[6] ), .A(\REGF/pbmemcnt1/sub_48/carry[6] 
        ), .B(\REGF/pbmemcnt1/down_data[6] ) );
    snl_or02x1 \REGF/pbmemcnt1/sub_48/U13  ( .Z(
        \REGF/pbmemcnt1/sub_48/carry[4] ), .A(\REGF/pbmemcnt1/down_data[3] ), 
        .B(\REGF/pbmemcnt1/sub_48/carry[3] ) );
    snl_or02x1 \REGF/pbmemcnt1/sub_48/U9  ( .Z(
        \REGF/pbmemcnt1/sub_48/carry[6] ), .A(\REGF/pbmemcnt1/down_data[5] ), 
        .B(\REGF/pbmemcnt1/sub_48/carry[5] ) );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U12  ( .ZN(
        \REGF/pbmemcnt1/down_data274[4] ), .A(\REGF/pbmemcnt1/sub_48/carry[4] 
        ), .B(\REGF/pbmemcnt1/down_data[4] ) );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U10  ( .ZN(
        \REGF/pbmemcnt1/down_data274[5] ), .A(\REGF/pbmemcnt1/sub_48/carry[5] 
        ), .B(\REGF/pbmemcnt1/down_data[5] ) );
    snl_or02x1 \REGF/pbmemcnt1/sub_48/U15  ( .Z(
        \REGF/pbmemcnt1/sub_48/carry[3] ), .A(\REGF/pbmemcnt1/down_data[2] ), 
        .B(\REGF/pbmemcnt1/sub_48/carry[2] ) );
    snl_or02x1 \REGF/pbmemcnt1/sub_48/U17  ( .Z(
        \REGF/pbmemcnt1/sub_48/carry[2] ), .A(\REGF/pbmemcnt1/down_data[1] ), 
        .B(\REGF/pbmemcnt1/down_data[0] ) );
    snl_or02x1 \REGF/pbmemcnt1/sub_48/U11  ( .Z(
        \REGF/pbmemcnt1/sub_48/carry[5] ), .A(\REGF/pbmemcnt1/down_data[4] ), 
        .B(\REGF/pbmemcnt1/sub_48/carry[4] ) );
    snl_invx05 \REGF/pbmemcnt1/sub_48/U19  ( .ZN(
        \REGF/pbmemcnt1/down_data274[0] ), .A(\REGF/pbmemcnt1/down_data[0] )
         );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U16  ( .ZN(
        \REGF/pbmemcnt1/down_data274[2] ), .A(\REGF/pbmemcnt1/sub_48/carry[2] 
        ), .B(\REGF/pbmemcnt1/down_data[2] ) );
    snl_xnor2x0 \REGF/pbmemcnt1/sub_48/U18  ( .ZN(
        \REGF/pbmemcnt1/down_data274[1] ), .A(\REGF/pbmemcnt1/down_data[0] ), 
        .B(\REGF/pbmemcnt1/down_data[1] ) );
    snl_invx05 \REG_2/SATIME/add_187/U5  ( .ZN(\REG_2/SATIME/count145[0] ), 
        .A(\REG_2/SATIME/count[0] ) );
    snl_xor2x0 \REG_2/SATIME/add_187/U6  ( .Z(\REG_2/SATIME/count145[20] ), 
        .A(\REG_2/SATIME/count[20] ), .B(\REG_2/SATIME/add_187/carry[20] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_10  ( .S(
        \REG_2/SATIME/count145[10] ), .CO(\REG_2/SATIME/add_187/carry[11] ), 
        .A(\REG_2/SATIME/count[10] ), .B(\REG_2/SATIME/add_187/carry[10] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_19  ( .S(
        \REG_2/SATIME/count145[19] ), .CO(\REG_2/SATIME/add_187/carry[20] ), 
        .A(\REG_2/SATIME/count[19] ), .B(\REG_2/SATIME/add_187/carry[19] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_3  ( .S(\REG_2/SATIME/count145[3] ), 
        .CO(\REG_2/SATIME/add_187/carry[4] ), .A(\REG_2/SATIME/count[3] ), .B(
        \REG_2/SATIME/add_187/carry[3] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_4  ( .S(\REG_2/SATIME/count145[4] ), 
        .CO(\REG_2/SATIME/add_187/carry[5] ), .A(\REG_2/SATIME/count[4] ), .B(
        \REG_2/SATIME/add_187/carry[4] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_17  ( .S(
        \REG_2/SATIME/count145[17] ), .CO(\REG_2/SATIME/add_187/carry[18] ), 
        .A(\REG_2/SATIME/count[17] ), .B(\REG_2/SATIME/add_187/carry[17] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_2  ( .S(\REG_2/SATIME/count145[2] ), 
        .CO(\REG_2/SATIME/add_187/carry[3] ), .A(\REG_2/SATIME/count[2] ), .B(
        \REG_2/SATIME/add_187/carry[2] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_5  ( .S(\REG_2/SATIME/count145[5] ), 
        .CO(\REG_2/SATIME/add_187/carry[6] ), .A(\REG_2/SATIME/count[5] ), .B(
        \REG_2/SATIME/add_187/carry[5] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_11  ( .S(
        \REG_2/SATIME/count145[11] ), .CO(\REG_2/SATIME/add_187/carry[12] ), 
        .A(\REG_2/SATIME/count[11] ), .B(\REG_2/SATIME/add_187/carry[11] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_16  ( .S(
        \REG_2/SATIME/count145[16] ), .CO(\REG_2/SATIME/add_187/carry[17] ), 
        .A(\REG_2/SATIME/count[16] ), .B(\REG_2/SATIME/add_187/carry[16] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_7  ( .S(\REG_2/SATIME/count145[7] ), 
        .CO(\REG_2/SATIME/add_187/carry[8] ), .A(\REG_2/SATIME/count[7] ), .B(
        \REG_2/SATIME/add_187/carry[7] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_13  ( .S(
        \REG_2/SATIME/count145[13] ), .CO(\REG_2/SATIME/add_187/carry[14] ), 
        .A(\REG_2/SATIME/count[13] ), .B(\REG_2/SATIME/add_187/carry[13] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_18  ( .S(
        \REG_2/SATIME/count145[18] ), .CO(\REG_2/SATIME/add_187/carry[19] ), 
        .A(\REG_2/SATIME/count[18] ), .B(\REG_2/SATIME/add_187/carry[18] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_1  ( .S(\REG_2/SATIME/count145[1] ), 
        .CO(\REG_2/SATIME/add_187/carry[2] ), .A(\REG_2/SATIME/count[1] ), .B(
        \REG_2/SATIME/count[0] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_9  ( .S(\REG_2/SATIME/count145[9] ), 
        .CO(\REG_2/SATIME/add_187/carry[10] ), .A(\REG_2/SATIME/count[9] ), 
        .B(\REG_2/SATIME/add_187/carry[9] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_14  ( .S(
        \REG_2/SATIME/count145[14] ), .CO(\REG_2/SATIME/add_187/carry[15] ), 
        .A(\REG_2/SATIME/count[14] ), .B(\REG_2/SATIME/add_187/carry[14] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_6  ( .S(\REG_2/SATIME/count145[6] ), 
        .CO(\REG_2/SATIME/add_187/carry[7] ), .A(\REG_2/SATIME/count[6] ), .B(
        \REG_2/SATIME/add_187/carry[6] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_8  ( .S(\REG_2/SATIME/count145[8] ), 
        .CO(\REG_2/SATIME/add_187/carry[9] ), .A(\REG_2/SATIME/count[8] ), .B(
        \REG_2/SATIME/add_187/carry[8] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_15  ( .S(
        \REG_2/SATIME/count145[15] ), .CO(\REG_2/SATIME/add_187/carry[16] ), 
        .A(\REG_2/SATIME/count[15] ), .B(\REG_2/SATIME/add_187/carry[15] ) );
    snl_add05x1 \REG_2/SATIME/add_187/U1_1_12  ( .S(
        \REG_2/SATIME/count145[12] ), .CO(\REG_2/SATIME/add_187/carry[13] ), 
        .A(\REG_2/SATIME/count[12] ), .B(\REG_2/SATIME/add_187/carry[12] ) );
    snl_ao012x1 \SAEXE/RFIO/phcont4_1/U28  ( .Z(
        \SAEXE/RFIO/phcont4_1/count52[0] ), .A(\SAEXE/RFIO/phcont4_1/ncnt[0] ), 
        .B(\SAEXE/RFIO/phcont4_1/n84 ), .C(\SAEXE/RFIO/cntloadh ) );
    snl_invx05 \SAEXE/RFIO/phcont4_1/U33  ( .ZN(\SAEXE/RFIO/phcont4_1/n86 ), 
        .A(\SAEXE/RFIO/phcont4_1/count[0] ) );
    snl_nand13x1 \SAEXE/RFIO/phcont4_1/U26  ( .ZN(\SAEXE/RFIO/phcont4_1/n_42 ), 
        .A(\SAEXE/RFIO/cnt4dech ), .B(\SAEXE/RFIO/phcont4_1/n83 ), .C(
        \SAEXE/RFIO/phcont4_1/n84 ) );
    snl_invx05 \SAEXE/RFIO/phcont4_1/U34  ( .ZN(\SAEXE/RFIO/phcont4_1/n87 ), 
        .A(\SAEXE/RFIO/phcont4_1/count[1] ) );
    snl_sffqensnx2 \SAEXE/RFIO/phcont4_1/count_reg[0]  ( .Q(
        \SAEXE/RFIO/phcont4_1/count[0] ), .D(1'b0), .EN(1'b1), .SN(n10735), 
        .SD(\SAEXE/RFIO/phcont4_1/count52[0] ), .SE(
        \SAEXE/RFIO/phcont4_1/n_42 ), .CP(SCLK) );
    snl_nand13x1 \SAEXE/RFIO/phcont4_1/U27  ( .ZN(
        \SAEXE/RFIO/phcont4_1/count52[1] ), .A(\SAEXE/RFIO/phcont4_1/ncnt[1] ), 
        .B(\SAEXE/RFIO/phcont4_1/n83 ), .C(\SAEXE/RFIO/phcont4_1/n84 ) );
    snl_invx05 \SAEXE/RFIO/phcont4_1/U35  ( .ZN(\SAEXE/RFIO/phcont4_1/n83 ), 
        .A(\SAEXE/RFIO/cntloadh ) );
    snl_nor02x1 \SAEXE/RFIO/phcont4_1/U29  ( .ZN(\SAEXE/RFIO/cnt4out[3] ), .A(
        \SAEXE/RFIO/phcont4_1/n86 ), .B(\SAEXE/RFIO/phcont4_1/n87 ) );
    snl_nor02x1 \SAEXE/RFIO/phcont4_1/U30  ( .ZN(\SAEXE/RFIO/cnt4out[2] ), .A(
        \SAEXE/RFIO/phcont4_1/count[0] ), .B(\SAEXE/RFIO/phcont4_1/n87 ) );
    snl_nor02x1 \SAEXE/RFIO/phcont4_1/U32  ( .ZN(\SAEXE/RFIO/cnt4out[0] ), .A(
        \SAEXE/RFIO/phcont4_1/count[1] ), .B(\SAEXE/RFIO/phcont4_1/count[0] )
         );
    snl_nor02x1 \SAEXE/RFIO/phcont4_1/U31  ( .ZN(\SAEXE/RFIO/cnt4out[1] ), .A(
        \SAEXE/RFIO/phcont4_1/count[1] ), .B(\SAEXE/RFIO/phcont4_1/n86 ) );
    snl_invx05 \SAEXE/RFIO/phcont4_1/U36  ( .ZN(\SAEXE/RFIO/phcont4_1/n84 ), 
        .A(\SAEXE/RFIO/reloadh ) );
    snl_sffqensnx2 \SAEXE/RFIO/phcont4_1/count_reg[1]  ( .Q(
        \SAEXE/RFIO/phcont4_1/count[1] ), .D(1'b0), .EN(1'b1), .SN(n10735), 
        .SD(\SAEXE/RFIO/phcont4_1/count52[1] ), .SE(
        \SAEXE/RFIO/phcont4_1/n_42 ), .CP(SCLK) );
    snl_and23x0 \SAEXE/RFIO/RIN1/U69  ( .Z(\SAEXE/RFIO/srcadr1_h ), .A(
        pktrscendh), .B(\SAEXE/RFIO/RIN1/n165 ), .C(\SAEXE/RFIO/rfio1h ) );
    snl_ao1b13x1 \SAEXE/RFIO/RIN1/U73  ( .Z(\SAEXE/RFIO/RIN1/nfst[0] ), .A(
        \SAEXE/rf_srcadr2_h ), .B(\SAEXE/RFIO/RIN1/n171 ), .C(
        \SAEXE/RFIO/RIN1/n172 ), .D(\SAEXE/RFIO/RIN1/n167 ), .E(
        \SAEXE/RFIO/ri1_trscdech ) );
    snl_invx05 \SAEXE/RFIO/RIN1/U74  ( .ZN(\SAEXE/RFIO/RIN1/n165 ), .A(
        \SAEXE/RFIO/RIN1/fst[1] ) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U83  ( .ZN(\SAEXE/RFIO/RIN1/n169 ), .A(
        pgadrovfh), .B(\SAEXE/RFIO/RIN1/fst[2] ) );
    snl_invx05 \SAEXE/RFIO/RIN1/U84  ( .ZN(\SAEXE/RFIO/phadrovfh ), .A(
        \SAEXE/RFIO/RIN1/n169 ) );
    snl_invx05 \SAEXE/RFIO/RIN1/U75  ( .ZN(\SAEXE/RFIO/RIN1/n171 ), .A(
        \SAEXE/RFIO/RIN1/fst[2] ) );
    snl_nor04x0 \SAEXE/RFIO/RIN1/U82  ( .ZN(\SAEXE/RFIO/ri1_trscdech ), .A(
        \SAEXE/RFIO/RIN1/n166 ), .B(\SAEXE/RFIO/RIN1/n165 ), .C(pktrscendh), 
        .D(\SAEXE/RFIO/rfin2h ) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U90  ( .ZN(\SAEXE/RFIO/RIN1/n176 ), .A(
        \SAEXE/RFIO/RIN1/n172 ), .B(\SAEXE/RFIO/RIN1/n171 ) );
    snl_oai012x1 \SAEXE/RFIO/RIN1/U70  ( .ZN(\SAEXE/RFIO/phrfin1sah ), .A(
        \SAEXE/RFIO/rfin1tpenh ), .B(\SAEXE/RFIO/RIN1/n166 ), .C(
        \SAEXE/RFIO/RIN1/n167 ) );
    snl_and34x0 \SAEXE/RFIO/RIN1/U72  ( .Z(\SAEXE/RFIO/RIN1/nfst[2] ), .A(
        \SAEXE/RFIO/RIN1/fst[2] ), .B(ph_lberr), .C(\SAEXE/RFIO/RIN1/n170 ), 
        .D(ph_lbend) );
    snl_oa012x1 \SAEXE/RFIO/RIN1/U85  ( .Z(\SAEXE/RFIO/rfin1tpenh ), .A(
        pktrscendh), .B(\SAEXE/RFIO/rfin2h ), .C(\SAEXE/RFIO/RIN1/fst[1] ) );
    snl_ffqrnx1 \SAEXE/RFIO/RIN1/fst_reg[1]  ( .Q(\SAEXE/RFIO/RIN1/fst[1] ), 
        .D(\SAEXE/RFIO/RIN1/nfst[1] ), .RN(n10735), .CP(SCLK) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U71  ( .ZN(\SAEXE/RFIO/phrefendh ), .A(
        \SAEXE/RFIO/RIN1/n168 ), .B(\SAEXE/RFIO/RIN1/n169 ) );
    snl_nand12x1 \SAEXE/RFIO/RIN1/U76  ( .ZN(\SAEXE/RFIO/RIN1/n166 ), .A(
        pgadrovfh), .B(\SAEXE/RFIO/RIN1/fst[2] ) );
    snl_nor02x1 \SAEXE/RFIO/RIN1/U77  ( .ZN(\SAEXE/RFIO/RIN1/n170 ), .A(
        \SAEXE/RFIO/RIN1/fst[1] ), .B(\SAEXE/rf_srcadr2_h ) );
    snl_muxi21x1 \SAEXE/RFIO/RIN1/U79  ( .ZN(\SAEXE/relbwrh ), .A(
        \SAEXE/RFIO/RIN1/n173 ), .B(\SAEXE/RFIO/RIN1/n174 ), .S(
        \SAEXE/rf_srcadr2_h ) );
    snl_ffqrnx1 \SAEXE/RFIO/RIN1/fst_reg[0]  ( .Q(\SAEXE/rf_srcadr2_h ), .D(
        \SAEXE/RFIO/RIN1/nfst[0] ), .RN(n10735), .CP(SCLK) );
    snl_nor02x1 \SAEXE/RFIO/RIN1/U80  ( .ZN(\SAEXE/RFIO/RIN1/n175 ), .A(
        \SAEXE/RFIO/RIN1/n170 ), .B(\SAEXE/RFIO/RIN1/n172 ) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U87  ( .ZN(\SAEXE/RFIO/RIN1/n174 ), .A(
        \SAEXE/RFIO/RIN1/fst[2] ), .B(\SAEXE/RFIO/RIN1/n165 ) );
    snl_aoi022x1 \SAEXE/RFIO/RIN1/U89  ( .ZN(\SAEXE/RFIO/RIN1/n168 ), .A(
        \SAEXE/RFIO/rfin1tpenh ), .B(\SAEXE/RFIO/RIN1/fst[2] ), .C(
        \SAEXE/RFIO/RIN1/n175 ), .D(\SAEXE/RFIO/RIN1/n171 ) );
    snl_ffqrnx1 \SAEXE/RFIO/RIN1/fst_reg[2]  ( .Q(\SAEXE/RFIO/RIN1/fst[2] ), 
        .D(\SAEXE/RFIO/RIN1/nfst[2] ), .RN(n10735), .CP(SCLK) );
    snl_aoi022x1 \SAEXE/RFIO/RIN1/U81  ( .ZN(\SAEXE/RFIO/RIN1/nfst[1] ), .A(
        \SAEXE/RFIO/RIN1/n176 ), .B(\SAEXE/RFIO/RIN1/fst[1] ), .C(
        \SAEXE/RFIO/RIN1/n166 ), .D(\SAEXE/RFIO/RIN1/n165 ) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U88  ( .ZN(\SAEXE/RFIO/RIN1/n173 ), .A(
        \SAEXE/RFIO/RIN1/fst[1] ), .B(\SAEXE/RFIO/RIN1/n171 ) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U78  ( .ZN(\SAEXE/RFIO/RIN1/n172 ), .A(
        ph_lbend), .B(ph_lberr) );
    snl_nand02x1 \SAEXE/RFIO/RIN1/U86  ( .ZN(\SAEXE/RFIO/RIN1/n167 ), .A(
        \SAEXE/RFIO/phrfin1h ), .B(\SAEXE/RFIO/RIN1/n170 ) );
    snl_ao012x1 \SADR/MAINSADR/addidxof/U6  ( .Z(
        \SADR/MAINSADR/addidxof/cin_stg[2] ), .A(
        \SADR/MAINSADR/addidxof/gp_out[2] ), .B(
        \SADR/MAINSADR/addidxof/cin_stg[1] ), .C(
        \SADR/MAINSADR/addidxof/gg_out[2] ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/U8  ( .ZN(
        \SADR/MAINSADR/addidxof/n8632 ), .A(\SADR/MAINSADR/addidxof/gp_out[3] 
        ), .B(\SADR/MAINSADR/addidxof/cin_stg[2] ), .C(
        \SADR/MAINSADR/addidxof/gg_out[3] ) );
    snl_ao012x1 \SADR/MAINSADR/addidxof/U7  ( .Z(
        \SADR/MAINSADR/addidxof/cin_stg[1] ), .A(
        \SADR/MAINSADR/addidxof/gp_out[1] ), .B(
        \SADR/MAINSADR/addidxof/gg_out[0] ), .C(
        \SADR/MAINSADR/addidxof/gg_out[1] ) );
    snl_xnor2x0 \SADR/MAINSADR/addidxof/U9  ( .ZN(
        \SADR/MAINSADR/ovf_addindoff ), .A(\SADR/MAINSADR/addidxof/c_last ), 
        .B(\SADR/MAINSADR/addidxof/n8632 ) );
    snl_and02x1 \SADR/MAINSADR/addsegoff/U6  ( .Z(
        \SADR/MAINSADR/addsegoff/n8497 ), .A(\SADR/MAINSADR/addsegoff/n8498 ), 
        .B(\SADR/segbase[16] ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/U14  ( .Z(\SADR/sadr[26] ), .A(
        \SADR/segbase[16] ), .B(\SADR/MAINSADR/addsegoff/n8498 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/U7  ( .ZN(
        \SADR/MAINSADR/addsegoff/n8499 ), .A(\SADR/MAINSADR/addsegoff/n8500 ), 
        .B(\SADR/MAINSADR/addsegoff/n8501 ) );
    snl_xnor2x0 \SADR/MAINSADR/addsegoff/U8  ( .ZN(\SADR/sadr[22] ), .A(
        \SADR/segbase[12] ), .B(\SADR/MAINSADR/addsegoff/n8502 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/U13  ( .Z(\SADR/sadr[27] ), .A(
        \SADR/MAINSADR/addsegoff/n8497 ), .B(\SADR/segbase[17] ) );
    snl_and12x1 \SADR/MAINSADR/addsegoff/U9  ( .Z(
        \SADR/MAINSADR/addsegoff/n8503 ), .A(\SADR/MAINSADR/addsegoff/n8502 ), 
        .B(\SADR/segbase[12] ) );
    snl_and23x0 \SADR/MAINSADR/addsegoff/U12  ( .Z(
        \SADR/MAINSADR/addsegoff/n8498 ), .A(\SADR/MAINSADR/addsegoff/n8501 ), 
        .B(\SADR/MAINSADR/addsegoff/n8500 ), .C(\SADR/segbase[15] ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/U10  ( .ZN(
        \SADR/MAINSADR/addsegoff/n8500 ), .A(\SADR/segbase[13] ), .B(
        \SADR/MAINSADR/addsegoff/n8503 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/U15  ( .Z(\SADR/sadr[25] ), .A(
        \SADR/segbase[15] ), .B(\SADR/MAINSADR/addsegoff/n8499 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/U17  ( .Z(\SADR/sadr[23] ), .A(
        \SADR/segbase[13] ), .B(\SADR/MAINSADR/addsegoff/n8503 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/U11  ( .ZN(
        \SADR/MAINSADR/addsegoff/n8501 ), .A(\SADR/segbase[14] ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/U18  ( .ZN(
        \SADR/MAINSADR/addsegoff/n8502 ), .A(
        \SADR/MAINSADR/addsegoff/gp_out[1] ), .B(
        \SADR/MAINSADR/addsegoff/gg_out[0] ), .C(
        \SADR/MAINSADR/addsegoff/gg_out[1] ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/U16  ( .Z(\SADR/sadr[24] ), .A(
        \SADR/MAINSADR/addsegoff/n8501 ), .B(\SADR/MAINSADR/addsegoff/n8500 )
         );
    snl_and02x1 \SADR/MAINSADR/adrinc1/U6  ( .Z(
        \SADR/MAINSADR/adrinc1/gg_out[4] ), .A(
        \SADR/MAINSADR/adrinc1/gp_out[4] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[3] ) );
    snl_and02x1 \SADR/MAINSADR/adrinc1/U8  ( .Z(
        \SADR/MAINSADR/adrinc1/gg_out[2] ), .A(
        \SADR/MAINSADR/adrinc1/gp_out[2] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[1] ) );
    snl_and02x1 \SADR/MAINSADR/adrinc1/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/gg_out[1] ), .A(
        \SADR/MAINSADR/adrinc1/gp_out[0] ), .B(
        \SADR/MAINSADR/adrinc1/gp_out[1] ) );
    snl_and02x1 \SADR/MAINSADR/adrinc1/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/gg_out[3] ), .A(
        \SADR/MAINSADR/adrinc1/gp_out[3] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[2] ) );
    snl_oa012x1 \SADR/MAINSADR/adrcmp1/U8  ( .Z(\SADR/MAINSADR/adrcmp1/n8405 ), 
        .A(\SADR/MAINSADR/adrcmp1/geq[0] ), .B(\SADR/MAINSADR/adrcmp1/ggfl[0] 
        ), .C(\SADR/MAINSADR/adrcmp1/geq[1] ) );
    snl_nand12x1 \SADR/MAINSADR/adrcmp1/U7  ( .ZN(\SADR/MAINSADR/cmpflg ), .A(
        \SADR/MAINSADR/adrcmp1/ggfl[3] ), .B(\SADR/MAINSADR/adrcmp1/n8404 ) );
    snl_oa012x1 \SADR/MAINSADR/adrcmp1/U9  ( .Z(\SADR/MAINSADR/adrcmp1/n8406 ), 
        .A(\SADR/MAINSADR/adrcmp1/n8405 ), .B(\SADR/MAINSADR/adrcmp1/ggfl[1] ), 
        .C(\SADR/MAINSADR/adrcmp1/geq[2] ) );
    snl_oai012x1 \SADR/MAINSADR/adrcmp1/U10  ( .ZN(
        \SADR/MAINSADR/adrcmp1/n8404 ), .A(\SADR/MAINSADR/adrcmp1/n8406 ), .B(
        \SADR/MAINSADR/adrcmp1/ggfl[2] ), .C(\SADR/MAINSADR/adrcmp1/geq[3] )
         );
    snl_or02x1 \SADR/MAINSADR/adrdec1/U6  ( .Z(
        \SADR/MAINSADR/adrdec1/gcarry[1] ), .A(
        \SADR/MAINSADR/adrdec1/gg_out[0] ), .B(
        \SADR/MAINSADR/adrdec1/gg_out[1] ) );
    snl_or02x1 \SADR/MAINSADR/adrdec1/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/gcarry[2] ), .A(
        \SADR/MAINSADR/adrdec1/gg_out[2] ), .B(
        \SADR/MAINSADR/adrdec1/gcarry[1] ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/U9  ( .ZN(\SADR/MAINSADR/adrdec1/n8347 
        ), .A(\SADR/MAINSADR/adrdec1/gg_out[3] ), .B(
        \SADR/MAINSADR/adrdec1/gcarry[2] ) );
    snl_nand12x1 \SADR/MAINSADR/adrdec1/U7  ( .ZN(
        \SADR/MAINSADR/adrdec1/gcarry[4] ), .A(
        \SADR/MAINSADR/adrdec1/gg_out[4] ), .B(\SADR/MAINSADR/adrdec1/n8347 )
         );
    snl_invx05 \SADR/MAINSADR/adrdec1/U10  ( .ZN(
        \SADR/MAINSADR/adrdec1/gcarry[3] ), .A(\SADR/MAINSADR/adrdec1/n8347 )
         );
    snl_and02x1 \SADR/MAINSADR/adrinc2/U6  ( .Z(
        \SADR/MAINSADR/adrinc2/gg_out[4] ), .A(
        \SADR/MAINSADR/adrinc2/gp_out[4] ), .B(
        \SADR/MAINSADR/adrinc2/gg_out[3] ) );
    snl_and02x1 \SADR/MAINSADR/adrinc2/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/gg_out[1] ), .A(
        \SADR/MAINSADR/adrinc2/gp_out[0] ), .B(
        \SADR/MAINSADR/adrinc2/gp_out[1] ) );
    snl_and02x1 \SADR/MAINSADR/adrinc2/U8  ( .Z(
        \SADR/MAINSADR/adrinc2/gg_out[2] ), .A(
        \SADR/MAINSADR/adrinc2/gp_out[2] ), .B(
        \SADR/MAINSADR/adrinc2/gg_out[1] ) );
    snl_and02x1 \SADR/MAINSADR/adrinc2/U9  ( .Z(
        \SADR/MAINSADR/adrinc2/gg_out[3] ), .A(
        \SADR/MAINSADR/adrinc2/gp_out[3] ), .B(
        \SADR/MAINSADR/adrinc2/gg_out[2] ) );
    snl_or02x1 \SADR/MAINSADR/adrdec2/U6  ( .Z(
        \SADR/MAINSADR/adrdec2/gcarry[1] ), .A(
        \SADR/MAINSADR/adrdec2/gg_out[0] ), .B(
        \SADR/MAINSADR/adrdec2/gg_out[1] ) );
    snl_or02x1 \SADR/MAINSADR/adrdec2/U8  ( .Z(
        \SADR/MAINSADR/adrdec2/gcarry[2] ), .A(
        \SADR/MAINSADR/adrdec2/gg_out[2] ), .B(
        \SADR/MAINSADR/adrdec2/gcarry[1] ) );
    snl_nand12x1 \SADR/MAINSADR/adrdec2/U7  ( .ZN(
        \SADR/MAINSADR/adrdec2/gcarry[4] ), .A(
        \SADR/MAINSADR/adrdec2/gg_out[4] ), .B(\SADR/MAINSADR/adrdec2/n8299 )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/U9  ( .ZN(\SADR/MAINSADR/adrdec2/n8299 
        ), .A(\SADR/MAINSADR/adrdec2/gg_out[3] ), .B(
        \SADR/MAINSADR/adrdec2/gcarry[2] ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/U10  ( .ZN(
        \SADR/MAINSADR/adrdec2/gcarry[3] ), .A(\SADR/MAINSADR/adrdec2/n8299 )
         );
    snl_and02x1 \REGF/pbmemff21/pbinc19k_1/U6  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gg_out[3] ), .A(
        \REGF/pbmemff21/pbinc19k_1/gp_out[3] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gg_out[2] ) );
    snl_and02x1 \REGF/pbmemff21/pbinc19k_1/U7  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gg_out[1] ), .A(
        \REGF/pbmemff21/pbinc19k_1/gp_out[1] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gp_out[0] ) );
    snl_and02x1 \REGF/pbmemff21/pbinc19k_1/U8  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gg_out[2] ), .A(
        \REGF/pbmemff21/pbinc19k_1/gp_out[2] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gg_out[1] ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x/U6  ( .Z(\SADR/ADDIDX/add_w_x/cin_stg[2] 
        ), .A(\SADR/ADDIDX/add_w_x/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_x/cin_stg[1] ), .C(\SADR/ADDIDX/add_w_x/gg_out[2] )
         );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/U8  ( .ZN(\SADR/ADDIDX/add_w_x/n10655 ), 
        .A(\SADR/ADDIDX/add_w_x/gp_out[3] ), .B(
        \SADR/ADDIDX/add_w_x/cin_stg[2] ), .C(\SADR/ADDIDX/add_w_x/gg_out[3] )
         );
    snl_ao012x1 \SADR/ADDIDX/add_w_x/U7  ( .Z(\SADR/ADDIDX/add_w_x/cin_stg[1] 
        ), .A(\SADR/ADDIDX/add_w_x/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_x/gg_out[0] ), .C(\SADR/ADDIDX/add_w_x/gg_out[1] )
         );
    snl_xnor2x0 \SADR/ADDIDX/add_w_x/U9  ( .ZN(\SADR/pgovfwx ), .A(
        \SADR/ADDIDX/add_w_x/c_last ), .B(\SADR/ADDIDX/add_w_x/n10655 ) );
    snl_ao012x1 \SADR/ADDIDX/add_x_z/U6  ( .Z(\SADR/ADDIDX/add_x_z/cin_stg[2] 
        ), .A(\SADR/ADDIDX/add_x_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_x_z/cin_stg[1] ), .C(\SADR/ADDIDX/add_x_z/gg_out[2] )
         );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/U8  ( .ZN(\SADR/ADDIDX/add_x_z/n10526 ), 
        .A(\SADR/ADDIDX/add_x_z/gp_out[3] ), .B(
        \SADR/ADDIDX/add_x_z/cin_stg[2] ), .C(\SADR/ADDIDX/add_x_z/gg_out[3] )
         );
    snl_ao012x1 \SADR/ADDIDX/add_x_z/U7  ( .Z(\SADR/ADDIDX/add_x_z/cin_stg[1] 
        ), .A(\SADR/ADDIDX/add_x_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_x_z/gg_out[0] ), .C(\SADR/ADDIDX/add_x_z/gg_out[1] )
         );
    snl_xnor2x0 \SADR/ADDIDX/add_x_z/U9  ( .ZN(\SADR/pgovfxz ), .A(
        \SADR/ADDIDX/add_x_z/c_last ), .B(\SADR/ADDIDX/add_x_z/n10526 ) );
    snl_ao012x1 \SADR/ADDIDX/add_y_z/U6  ( .Z(\SADR/ADDIDX/add_y_z/cin_stg[2] 
        ), .A(\SADR/ADDIDX/add_y_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_y_z/cin_stg[1] ), .C(\SADR/ADDIDX/add_y_z/gg_out[2] )
         );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/U8  ( .ZN(\SADR/ADDIDX/add_y_z/n10397 ), 
        .A(\SADR/ADDIDX/add_y_z/gp_out[3] ), .B(
        \SADR/ADDIDX/add_y_z/cin_stg[2] ), .C(\SADR/ADDIDX/add_y_z/gg_out[3] )
         );
    snl_ao012x1 \SADR/ADDIDX/add_y_z/U7  ( .Z(\SADR/ADDIDX/add_y_z/cin_stg[1] 
        ), .A(\SADR/ADDIDX/add_y_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_y_z/gg_out[0] ), .C(\SADR/ADDIDX/add_y_z/gg_out[1] )
         );
    snl_xnor2x0 \SADR/ADDIDX/add_y_z/U9  ( .ZN(\SADR/pgovfyz ), .A(
        \SADR/ADDIDX/add_y_z/c_last ), .B(\SADR/ADDIDX/add_y_z/n10397 ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_y/U6  ( .Z(\SADR/ADDIDX/add_w_y/cin_stg[2] 
        ), .A(\SADR/ADDIDX/add_w_y/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_y/cin_stg[1] ), .C(\SADR/ADDIDX/add_w_y/gg_out[2] )
         );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/U8  ( .ZN(\SADR/ADDIDX/add_w_y/n10268 ), 
        .A(\SADR/ADDIDX/add_w_y/gp_out[3] ), .B(
        \SADR/ADDIDX/add_w_y/cin_stg[2] ), .C(\SADR/ADDIDX/add_w_y/gg_out[3] )
         );
    snl_ao012x1 \SADR/ADDIDX/add_w_y/U7  ( .Z(\SADR/ADDIDX/add_w_y/cin_stg[1] 
        ), .A(\SADR/ADDIDX/add_w_y/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_y/gg_out[0] ), .C(\SADR/ADDIDX/add_w_y/gg_out[1] )
         );
    snl_xnor2x0 \SADR/ADDIDX/add_w_y/U9  ( .ZN(\SADR/pgovfwy ), .A(
        \SADR/ADDIDX/add_w_y/c_last ), .B(\SADR/ADDIDX/add_w_y/n10268 ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x_y/U6  ( .Z(
        \SADR/ADDIDX/add_w_x_y/cin_stg[2] ), .A(
        \SADR/ADDIDX/add_w_x_y/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_x_y/cin_stg[1] ), .C(
        \SADR/ADDIDX/add_w_x_y/gg_out[2] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/n10139 ), .A(\SADR/ADDIDX/add_w_x_y/gp_out[3] ), 
        .B(\SADR/ADDIDX/add_w_x_y/cin_stg[2] ), .C(
        \SADR/ADDIDX/add_w_x_y/gg_out[3] ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x_y/U7  ( .Z(
        \SADR/ADDIDX/add_w_x_y/cin_stg[1] ), .A(
        \SADR/ADDIDX/add_w_x_y/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_x_y/gg_out[0] ), .C(
        \SADR/ADDIDX/add_w_x_y/gg_out[1] ) );
    snl_xnor2x0 \SADR/ADDIDX/add_w_x_y/U9  ( .ZN(\SADR/ADDIDX/pgovfwxyT ), .A(
        \SADR/ADDIDX/add_w_x_y/c_last ), .B(\SADR/ADDIDX/add_w_x_y/n10139 ) );
    snl_ao012x1 \SADR/ADDIDX/add_x_y_z/U6  ( .Z(
        \SADR/ADDIDX/add_x_y_z/cin_stg[2] ), .A(
        \SADR/ADDIDX/add_x_y_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_x_y_z/cin_stg[1] ), .C(
        \SADR/ADDIDX/add_x_y_z/gg_out[2] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/n10010 ), .A(\SADR/ADDIDX/add_x_y_z/gp_out[3] ), 
        .B(\SADR/ADDIDX/add_x_y_z/cin_stg[2] ), .C(
        \SADR/ADDIDX/add_x_y_z/gg_out[3] ) );
    snl_ao012x1 \SADR/ADDIDX/add_x_y_z/U7  ( .Z(
        \SADR/ADDIDX/add_x_y_z/cin_stg[1] ), .A(
        \SADR/ADDIDX/add_x_y_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_x_y_z/gg_out[0] ), .C(
        \SADR/ADDIDX/add_x_y_z/gg_out[1] ) );
    snl_xnor2x0 \SADR/ADDIDX/add_x_y_z/U9  ( .ZN(\SADR/ADDIDX/pgovfxyzT ), .A(
        \SADR/ADDIDX/add_x_y_z/c_last ), .B(\SADR/ADDIDX/add_x_y_z/n10010 ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_z/U6  ( .Z(\SADR/ADDIDX/add_w_z/cin_stg[2] 
        ), .A(\SADR/ADDIDX/add_w_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_z/cin_stg[1] ), .C(\SADR/ADDIDX/add_w_z/gg_out[2] )
         );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/U8  ( .ZN(\SADR/ADDIDX/add_w_z/n9881 ), 
        .A(\SADR/ADDIDX/add_w_z/gp_out[3] ), .B(
        \SADR/ADDIDX/add_w_z/cin_stg[2] ), .C(\SADR/ADDIDX/add_w_z/gg_out[3] )
         );
    snl_ao012x1 \SADR/ADDIDX/add_w_z/U7  ( .Z(\SADR/ADDIDX/add_w_z/cin_stg[1] 
        ), .A(\SADR/ADDIDX/add_w_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_z/gg_out[0] ), .C(\SADR/ADDIDX/add_w_z/gg_out[1] )
         );
    snl_xnor2x0 \SADR/ADDIDX/add_w_z/U9  ( .ZN(\SADR/pgovfwz ), .A(
        \SADR/ADDIDX/add_w_z/c_last ), .B(\SADR/ADDIDX/add_w_z/n9881 ) );
    snl_ao012x1 \SADR/ADDIDX/add_x_y/U6  ( .Z(\SADR/ADDIDX/add_x_y/cin_stg[2] 
        ), .A(\SADR/ADDIDX/add_x_y/gp_out[2] ), .B(
        \SADR/ADDIDX/add_x_y/cin_stg[1] ), .C(\SADR/ADDIDX/add_x_y/gg_out[2] )
         );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/U8  ( .ZN(\SADR/ADDIDX/add_x_y/n9752 ), 
        .A(\SADR/ADDIDX/add_x_y/gp_out[3] ), .B(
        \SADR/ADDIDX/add_x_y/cin_stg[2] ), .C(\SADR/ADDIDX/add_x_y/gg_out[3] )
         );
    snl_ao012x1 \SADR/ADDIDX/add_x_y/U7  ( .Z(\SADR/ADDIDX/add_x_y/cin_stg[1] 
        ), .A(\SADR/ADDIDX/add_x_y/gp_out[1] ), .B(
        \SADR/ADDIDX/add_x_y/gg_out[0] ), .C(\SADR/ADDIDX/add_x_y/gg_out[1] )
         );
    snl_xnor2x0 \SADR/ADDIDX/add_x_y/U9  ( .ZN(\SADR/pgovfxy ), .A(
        \SADR/ADDIDX/add_x_y/c_last ), .B(\SADR/ADDIDX/add_x_y/n9752 ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x_z/U6  ( .Z(
        \SADR/ADDIDX/add_w_x_z/cin_stg[2] ), .A(
        \SADR/ADDIDX/add_w_x_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_x_z/cin_stg[1] ), .C(
        \SADR/ADDIDX/add_w_x_z/gg_out[2] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/n9623 ), .A(\SADR/ADDIDX/add_w_x_z/gp_out[3] ), 
        .B(\SADR/ADDIDX/add_w_x_z/cin_stg[2] ), .C(
        \SADR/ADDIDX/add_w_x_z/gg_out[3] ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x_z/U7  ( .Z(
        \SADR/ADDIDX/add_w_x_z/cin_stg[1] ), .A(
        \SADR/ADDIDX/add_w_x_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_x_z/gg_out[0] ), .C(
        \SADR/ADDIDX/add_w_x_z/gg_out[1] ) );
    snl_xnor2x0 \SADR/ADDIDX/add_w_x_z/U9  ( .ZN(\SADR/ADDIDX/pgovfwxzT ), .A(
        \SADR/ADDIDX/add_w_x_z/c_last ), .B(\SADR/ADDIDX/add_w_x_z/n9623 ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_y_z/U6  ( .Z(
        \SADR/ADDIDX/add_w_y_z/cin_stg[2] ), .A(
        \SADR/ADDIDX/add_w_y_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_y_z/cin_stg[1] ), .C(
        \SADR/ADDIDX/add_w_y_z/gg_out[2] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/n9494 ), .A(\SADR/ADDIDX/add_w_y_z/gp_out[3] ), 
        .B(\SADR/ADDIDX/add_w_y_z/cin_stg[2] ), .C(
        \SADR/ADDIDX/add_w_y_z/gg_out[3] ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_y_z/U7  ( .Z(
        \SADR/ADDIDX/add_w_y_z/cin_stg[1] ), .A(
        \SADR/ADDIDX/add_w_y_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_y_z/gg_out[0] ), .C(
        \SADR/ADDIDX/add_w_y_z/gg_out[1] ) );
    snl_xnor2x0 \SADR/ADDIDX/add_w_y_z/U9  ( .ZN(\SADR/ADDIDX/pgovfwyzT ), .A(
        \SADR/ADDIDX/add_w_y_z/c_last ), .B(\SADR/ADDIDX/add_w_y_z/n9494 ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x_y_z/U6  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[2] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/gp_out[2] ), .B(
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[1] ), .C(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[2] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/n9365 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/gp_out[3] ), .B(
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[2] ), .C(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[3] ) );
    snl_ao012x1 \SADR/ADDIDX/add_w_x_y_z/U7  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[1] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/gp_out[1] ), .B(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[0] ), .C(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[1] ) );
    snl_xnor2x0 \SADR/ADDIDX/add_w_x_y_z/U9  ( .ZN(\SADR/ADDIDX/pgovfwxyzT ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y_z/n9365 ) );
    snl_oa012x1 \REGF/pbmemff41/phdec12_2/U6  ( .Z(pktrscovfh), .A(
        \REGF/pbmemff41/phdec12_2/n7080 ), .B(\pk_stdat[0] ), .C(
        \pk_stdat[11] ) );
    snl_or02x1 \REGF/pbmemff41/phdec12_2/U8  ( .Z(
        \REGF/pbmemff41/phdec12_2/gcarry[1] ), .A(
        \REGF/pbmemff41/phdec12_2/gg_out[0] ), .B(
        \REGF/pbmemff41/phdec12_2/gg_out[1] ) );
    snl_nor03x0 \REGF/pbmemff41/phdec12_2/U7  ( .ZN(pktrscendh), .A(
        \REGF/pbmemff41/phdec12_2/n7080 ), .B(\pk_stdat[11] ), .C(
        \pk_stdat[0] ) );
    snl_or08x1 \REGF/pbmemff41/phdec12_2/U9  ( .Z(
        \REGF/pbmemff41/phdec12_2/n7080 ), .A(\pk_stdat[1] ), .B(\pk_stdat[6] 
        ), .C(\pk_stdat[10] ), .D(\pk_stdat[9] ), .E(\pk_stdat[4] ), .F(
        \pk_stdat[2] ), .G(\pk_stdat[7] ), .H(\REGF/pbmemff41/phdec12_2/n7081 
        ) );
    snl_or03x1 \REGF/pbmemff41/phdec12_2/U10  ( .Z(
        \REGF/pbmemff41/phdec12_2/n7081 ), .A(\pk_stdat[8] ), .B(\pk_stdat[5] 
        ), .C(\pk_stdat[3] ) );
    snl_oa012x1 \REGF/pbmemff41/phdec12_1/U6  ( .Z(pktblcovfh), .A(
        \REGF/pbmemff41/phdec12_1/n7063 ), .B(\pk_stdat[12] ), .C(
        \REGF/RO_TRCO[27] ) );
    snl_or02x1 \REGF/pbmemff41/phdec12_1/U8  ( .Z(
        \REGF/pbmemff41/phdec12_1/gcarry[1] ), .A(
        \REGF/pbmemff41/phdec12_1/gg_out[0] ), .B(
        \REGF/pbmemff41/phdec12_1/gg_out[1] ) );
    snl_nor03x0 \REGF/pbmemff41/phdec12_1/U7  ( .ZN(pktblcendh), .A(
        \REGF/pbmemff41/phdec12_1/n7063 ), .B(\REGF/RO_TRCO[27] ), .C(
        \pk_stdat[12] ) );
    snl_or08x1 \REGF/pbmemff41/phdec12_1/U9  ( .Z(
        \REGF/pbmemff41/phdec12_1/n7063 ), .A(\pk_stdat[13] ), .B(
        \pk_stdat[18] ), .C(\REGF/RO_TRCO[26] ), .D(\REGF/RO_TRCO[25] ), .E(
        \pk_stdat[16] ), .F(\pk_stdat[14] ), .G(\pk_stdat[19] ), .H(
        \REGF/pbmemff41/phdec12_1/n7064 ) );
    snl_or03x1 \REGF/pbmemff41/phdec12_1/U10  ( .Z(
        \REGF/pbmemff41/phdec12_1/n7064 ), .A(\pk_stdat[20] ), .B(
        \pk_stdat[17] ), .C(\pk_stdat[15] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U191  ( .ZN(\MAIN/ENGIN/STEP_A/tmp2[0] ), 
        .A(\MAIN/ENGIN/STEP_A/n3546 ), .B(\MAIN/ENGIN/STEP_A/n3547 ) );
    snl_oai113x0 \MAIN/ENGIN/STEP_A/U198  ( .ZN(\MAIN/ENGIN/a_swctl_st ), .A(
        \MAIN/ENGIN/STEP_A/n3544 ), .B(\MAIN/exe_end ), .C(
        \MAIN/ENGIN/STEP_A/n3563 ), .D(\MAIN/ENGIN/STEP_A/n3564 ), .E(
        \MAIN/ENGIN/STEP_A/n3565 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_A/U204  ( .ZN(
        \MAIN/ENGIN/STEP_A/decode_stage272 ), .A(\MAIN/ENGIN/STEP_A/n3567 ), 
        .B(\MAIN/ENGIN/STEP_A/tmp2[2] ), .C(\MAIN/ENGIN/STEP_A/n3548 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_A/U223  ( .ZN(\MAIN/ENGIN/STEP_A/n3580 ), 
        .A(\MAIN/ENGIN/STEP_A/cst[0] ), .B(\MAIN/ENGIN/STEP_A/n3571 ), .C(
        \MAIN/ENGIN/STEP_A/n3577 ) );
    snl_aoi222x0 \MAIN/ENGIN/STEP_A/U238  ( .ZN(\MAIN/ENGIN/STEP_A/n3565 ), 
        .A(\MAIN/ENGIN/A_INIT_STAGE ), .B(\MAIN/ENGIN/STEP_A/n3578 ), .C(
        \MAIN/ENGIN/STEP_A/n3577 ), .D(\MAIN/ENGIN/STEP_A/n3576 ), .E(
        \MAIN/ENGIN/STEP_A/n3587 ), .F(\MAIN/ENGIN/STEP_A/n3571 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_A/U256  ( .ZN(\MAIN/ENGIN/STEP_A/n3585 ), 
        .A(\MAIN/ENGIN/STEP_A/n3557 ), .B(\MAIN/ENGIN/STEP_A/n3582 ), .C(
        \MAIN/ENGIN/STEP_A/n3575 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U196  ( .ZN(\MAIN/ENGIN/a_decctl_st ), .A(
        \MAIN/ENGIN/STEP_A/n3561 ), .B(\MAIN/ENGIN/STEP_A/n3562 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U211  ( .ZN(\MAIN/ENGIN/STEP_A/n3563 ), 
        .A(\MAIN/ENGIN/STEP_A/cst[1] ), .B(\MAIN/ENGIN/STEP_A/cst[0] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U216  ( .ZN(\MAIN/ENGIN/STEP_A/n3579 ), 
        .A(\MAIN/ENGIN/STEP_A/n3577 ), .B(\MAIN/ENGIN/STEP_A/n3569 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_A/U231  ( .ZN(\MAIN/ENGIN/STEP_A/n3574 ), .A(
        \MAIN/ENGIN/STEP_A/cst[2] ), .B(\MAIN/ENGIN/STEP_A/cst[3] ), .C(
        \MAIN/ENGIN/STEP_A/n3568 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U244  ( .ZN(\MAIN/ENGIN/cf_st2_rst ), .A(
        \MAIN/ENGIN/STEP_A/n3581 ) );
    snl_aoi122x0 \MAIN/ENGIN/STEP_A/U236  ( .ZN(\MAIN/ENGIN/STEP_A/n3546 ), 
        .A(pk_pexe01_h), .B(\MAIN/ENGIN/STEP_A/n3585 ), .C(
        \MAIN/ENGIN/STEP_A/n3556 ), .D(\MAIN/ENGIN/STEP_A/n3586 ), .E(
        \MAIN/ENGIN/STEP_A/n3555 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U243  ( .ZN(step1_cf), .A(
        \MAIN/ENGIN/STEP_A/n3581 ), .B(pgperrh) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U258  ( .ZN(\MAIN/ENGIN/STEP_A/n3567 ), .A(
        \MAIN/ENGIN/STEP_A/tmp2[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U218  ( .ZN(\MAIN/ENGIN/STEP_A/n3560 ), .A(
        pk_pexe01_h) );
    snl_ao1b1b3x0 \MAIN/ENGIN/STEP_A/U251  ( .Z(\MAIN/ENGIN/STEP_A/n3553 ), 
        .A(\MAIN/ENGIN/STEP_A/n3588 ), .B(\MAIN/ENGIN/cf_start ), .C(
        \MAIN/excep_valid ), .D(\MAIN/ENGIN/STEP_A/n3568 ), .E(
        \MAIN/ENGIN/STEP_A/n3590 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U190  ( .ZN(\MAIN/ENGIN/a_d2_stage ), .A(
        \MAIN/ENGIN/STEP_A/n3544 ), .B(\MAIN/ENGIN/STEP_A/n3545 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_A/U197  ( .ZN(\MAIN/ENGIN/a_exectl_st ), .A(
        \MAIN/ENGIN/STEP_A/n3556 ), .B(\MAIN/ENGIN/STEP_A/n3544 ), .C(
        \MAIN/ENGIN/STEP_A/n3554 ) );
    snl_ao112x1 \MAIN/ENGIN/STEP_A/U203  ( .Z(\MAIN/ENGIN/b_dec_start ), .A(
        \MAIN/ENGIN/STEP_A/n3568 ), .B(\MAIN/ENGIN/STEP_A/n3569 ), .C(
        \MAIN/ENGIN/STEP_A/n3554 ), .D(\MAIN/ENGIN/STEP_A/cst[2] ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_A/U224  ( .ZN(\MAIN/ENGIN/STEP_A/n3581 ), 
        .A(\MAIN/ENGIN/a_cf_stage ), .B(\MAIN/ENGIN/STEP_A/n3556 ), .C(
        pgiaendp) );
    snl_aoi112x0 \MAIN/ENGIN/STEP_A/U199  ( .ZN(\MAIN/ENGIN/dec_st2_rst ), .A(
        \MAIN/ENGIN/STEP_A/n3556 ), .B(\MAIN/ENGIN/STEP_A/n3566 ), .C(
        \MAIN/ENGIN/STEP_A/n3563 ), .D(\MAIN/ENGIN/STEP_A/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U202  ( .ZN(ph_dec_ah), .A(
        \MAIN/ENGIN/a_dec_stage ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U210  ( .ZN(\MAIN/ENGIN/STEP_A/n3568 ), .A(
        \MAIN/ENGIN/STEP_A/cst[1] ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U242  ( .ZN(\MAIN/ENGIN/a_step_end ), .A(
        \MAIN/ENGIN/STEP_A/n3558 ) );
    snl_ao022x1 \MAIN/ENGIN/STEP_A/U259  ( .Z(\MAIN/ENGIN/STEP_A/n3589 ), .A(
        \MAIN/exe_end ), .B(\MAIN/ENGIN/STEP_A/cst[2] ), .C(
        \MAIN/ENGIN/STEP_A/n3583 ), .D(\MAIN/ENGIN/STEP_A/n3544 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_A/cst_reg[0]  ( .Q(\MAIN/ENGIN/STEP_A/cst[0] 
        ), .D(\MAIN/ENGIN/STEP_A/tmp2[0] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U237  ( .ZN(\MAIN/ENGIN/STEP_A/n3564 ), .A(
        \MAIN/ENGIN/STEP_A/n3574 ), .B(\MAIN/ENGIN/STEP_A/n3550 ) );
    snl_and34x0 \MAIN/ENGIN/STEP_A/U205  ( .Z(\MAIN/ENGIN/STEP_A/n3570 ), .A(
        \MAIN/ENGIN/STEP_A/cst[1] ), .B(\MAIN/ENGIN/STEP_A/cst[0] ), .C(
        \MAIN/ENGIN/STEP_A/n3571 ), .D(\MAIN/POL_STH ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U219  ( .ZN(\MAIN/ENGIN/STEP_A/n3556 ), .A(
        \MAIN/ENGIN/STEP_A/n3560 ), .B(\MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U225  ( .ZN(\MAIN/ENGIN/STEP_A/n3582 ), 
        .A(\MAIN/ENGIN/STEP_A/cst[2] ), .B(\MAIN/ENGIN/STEP_A/n3568 ) );
    snl_aoi012x1 \MAIN/ENGIN/STEP_A/U250  ( .ZN(\MAIN/ENGIN/STEP_A/n3590 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/cf_start ), .C(
        \MAIN/ENGIN/STEP_A/n3573 ) );
    snl_ao01b2x0 \MAIN/ENGIN/STEP_A/U222  ( .Z(\MAIN/ENGIN/STEP_A/n3555 ), .A(
        \MAIN/ENGIN/STEP_A/n3578 ), .B(\MAIN/ENGIN/STEP_A/n3579 ), .C(
        \MAIN/ENGIN/status_wr1 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U239  ( .ZN(\MAIN/ENGIN/A_INIT_STAGE ), .A(
        \MAIN/ENGIN/STEP_A/n3579 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U257  ( .ZN(\MAIN/ENGIN/STEP_A/n3584 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/STEP_A/n3557 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U217  ( .ZN(\MAIN/ENGIN/STEP_A/n3571 ), .A(
        \MAIN/ENGIN/STEP_A/cst[3] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U230  ( .ZN(\MAIN/ENGIN/STEP_A/n3554 ), .A(
        \MAIN/ENGIN/STEP_A/n3566 ), .B(\MAIN/ENGIN/STEP_A/n3563 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U245  ( .ZN(\MAIN/ENGIN/STEP_A/n3588 ), .A(
        \MAIN/ENGIN/STEP_A/n3556 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_A/cst_reg[2]  ( .Q(\MAIN/ENGIN/STEP_A/cst[2] 
        ), .D(\MAIN/ENGIN/STEP_A/tmp2[2] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_A/exec_stage_reg  ( .Q(\MAIN/a_exec_stage ), 
        .D(\MAIN/ENGIN/STEP_A/exec_stage278 ), .RN(\MAIN/ENGIN/n3591 ), .CP(
        SCLK) );
    snl_and34x0 \MAIN/ENGIN/STEP_A/U192  ( .Z(\MAIN/ENGIN/STEP_A/n3548 ), .A(
        \MAIN/ENGIN/STEP_A/n3550 ), .B(\MAIN/ENGIN/STEP_A/n3551 ), .C(step1_cf
        ), .D(\MAIN/ENGIN/STEP_A/n3549 ) );
    snl_aoi013x0 \MAIN/ENGIN/STEP_A/U207  ( .ZN(\MAIN/ENGIN/STEP_A/n3561 ), 
        .A(\MAIN/ENGIN/STEP_A/n3556 ), .B(\MAIN/ENGIN/STEP_A/n3573 ), .C(
        \MAIN/ENGIN/STEP_A/n3574 ), .D(step1_cf) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U220  ( .ZN(\MAIN/ENGIN/STEP_A/n3557 ), .A(
        \MAIN/ENGIN/cf_start ) );
    snl_oai233x0 \MAIN/ENGIN/STEP_A/U255  ( .ZN(\MAIN/ENGIN/STEP_A/n3586 ), 
        .A(\MAIN/ENGIN/STEP_A/n3571 ), .B(\MAIN/ENGIN/A_PED4_BR ), .C(
        \MAIN/ENGIN/STEP_A/n3573 ), .D(\MAIN/ENGIN/STEP_A/n3562 ), .E(
        \MAIN/ENGIN/STEP_A/cst[2] ), .F(\MAIN/ENGIN/STEP_A/n3568 ), .G(
        \MAIN/ENGIN/STEP_A/n3572 ), .H(\MAIN/ENGIN/STEP_A/n3580 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_A/cst_reg[3]  ( .Q(\MAIN/ENGIN/STEP_A/cst[3] 
        ), .D(\MAIN/ENGIN/STEP_A/nst[3] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_A/U193  ( .ZN(\MAIN/ENGIN/STEP_A/n3552 ), 
        .A(\MAIN/ENGIN/STEP_A/cst[2] ), .B(\MAIN/ENGIN/STEP_A/n3553 ), .C(
        \MAIN/ENGIN/STEP_A/n3554 ), .D(\MAIN/ENGIN/STEP_A/n3555 ) );
    snl_ao023x1 \MAIN/ENGIN/STEP_A/U194  ( .Z(\MAIN/ENGIN/STEP_A/nst[3] ), .A(
        \MAIN/ENGIN/STEP_A/n3556 ), .B(\MAIN/ENGIN/STEP_A/n3545 ), .C(
        \MAIN/ENGIN/STEP_A/cst[3] ), .D(\MAIN/ENGIN/cf_st2_rst ), .E(pgperrh)
         );
    snl_oai022x1 \MAIN/ENGIN/STEP_A/U195  ( .ZN(\MAIN/ENGIN/a_cfctl_st ), .A(
        \MAIN/ENGIN/STEP_A/n3557 ), .B(\MAIN/ENGIN/STEP_A/n3558 ), .C(
        \MAIN/ENGIN/STEP_A/n3559 ), .D(\MAIN/ENGIN/STEP_A/n3560 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U212  ( .ZN(\MAIN/ENGIN/STEP_A/n3566 ), .A(
        \MAIN/dec_end ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_A/U215  ( .ZN(\MAIN/ENGIN/STEP_A/n3578 ), 
        .A(\MAIN/ENGIN/STEP_A/n3557 ), .B(\MAIN/ENGIN/STEP_A/n3560 ), .C(
        \MAIN/POL_STH ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U229  ( .ZN(\MAIN/ENGIN/STEP_A/n3562 ), .A(
        \MAIN/ENGIN/dec_start ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_A/decode_stage_reg  ( .Q(
        \MAIN/ENGIN/a_dec_stage ), .D(\MAIN/ENGIN/STEP_A/decode_stage272 ), 
        .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK) );
    snl_nor03x0 \MAIN/ENGIN/STEP_A/U247  ( .ZN(\MAIN/ENGIN/STEP_A/n3550 ), .A(
        \MAIN/ENGIN/STEP_A/n3568 ), .B(pol_status), .C(
        \MAIN/ENGIN/STEP_A/n3544 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U232  ( .ZN(\MAIN/ENGIN/STEP_A/n3545 ), 
        .A(\MAIN/ENGIN/STEP_A/cst[1] ), .B(\MAIN/ENGIN/STEP_A/n3573 ) );
    snl_aoi123x0 \MAIN/ENGIN/STEP_A/U235  ( .ZN(\MAIN/ENGIN/STEP_A/n3547 ), 
        .A(\MAIN/ENGIN/STEP_A/cst[2] ), .B(\MAIN/ENGIN/STEP_A/cst[1] ), .C(
        pol_status), .D(\MAIN/ENGIN/STEP_A/sw_stage ), .E(
        \MAIN/ENGIN/STEP_A/n3584 ), .F(\MAIN/ENGIN/STEP_A/n3551 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U240  ( .ZN(\MAIN/ENGIN/a_cf_stage ), .A(
        \MAIN/ENGIN/STEP_A/n3580 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_A/U200  ( .ZN(
        \MAIN/ENGIN/STEP_A/exec_stage278 ), .A(\MAIN/ENGIN/STEP_A/n3567 ), .B(
        \MAIN/ENGIN/STEP_A/n3552 ), .C(\MAIN/ENGIN/STEP_A/n3548 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U209  ( .ZN(\MAIN/ENGIN/STEP_A/n3573 ), .A(
        \MAIN/ENGIN/STEP_A/cst[0] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U227  ( .ZN(\MAIN/ENGIN/STEP_A/d3_stage ), 
        .A(\MAIN/ENGIN/STEP_A/n3582 ), .B(\MAIN/ENGIN/STEP_A/cst[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U249  ( .ZN(\MAIN/ENGIN/STEP_A/n3569 ), .A(
        \MAIN/ENGIN/STEP_A/n3576 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U252  ( .ZN(\MAIN/ENGIN/STEP_A/tmp2[2] ), 
        .A(\MAIN/ENGIN/STEP_A/n3552 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_A/cst_reg[1]  ( .Q(\MAIN/ENGIN/STEP_A/cst[1] 
        ), .D(\MAIN/ENGIN/STEP_A/tmp2[1] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_invx05 \MAIN/ENGIN/STEP_A/U201  ( .ZN(ph_exe_ah), .A(
        \MAIN/a_exec_stage ) );
    snl_aoi0b12x0 \MAIN/ENGIN/STEP_A/U208  ( .ZN(\MAIN/ENGIN/STEP_A/n3559 ), 
        .A(\MAIN/ENGIN/STEP_A/d3_stage ), .B(\MAIN/ENGIN/cf_start ), .C(
        \MAIN/ENGIN/STEP_A/n3575 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U213  ( .ZN(\MAIN/ENGIN/STEP_A/n3576 ), 
        .A(\MAIN/ENGIN/STEP_A/n3571 ), .B(\MAIN/ENGIN/STEP_A/n3573 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U234  ( .ZN(\MAIN/ENGIN/STEP_A/n3583 ), .A(
        \MAIN/dec_end ), .B(\MAIN/ENGIN/STEP_A/n3556 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U241  ( .ZN(\MAIN/ENGIN/status_wr1 ), .A(
        \MAIN/ENGIN/STEP_A/n3571 ), .B(\MAIN/ENGIN/STEP_A/n3568 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U226  ( .ZN(\MAIN/ENGIN/STEP_A/sw_stage ), 
        .A(\MAIN/ENGIN/STEP_A/n3582 ), .B(\MAIN/ENGIN/STEP_A/n3573 ) );
    snl_and23x0 \MAIN/ENGIN/STEP_A/U206  ( .Z(\MAIN/ENGIN/STEP_A/n3572 ), .A(
        \MAIN/ENGIN/dec_start ), .B(pgperrh), .C(pgiaendp) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U248  ( .ZN(\MAIN/ENGIN/STEP_A/n3587 ), .A(
        \MAIN/ENGIN/STEP_A/n3582 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_A/U253  ( .ZN(\MAIN/ENGIN/STEP_A/n3549 ), 
        .A(\MAIN/ENGIN/STEP_A/n3570 ), .B(\MAIN/ENGIN/STEP_A/n3574 ), .C(
        \MAIN/ENGIN/STEP_A/n3556 ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U254  ( .ZN(\MAIN/ENGIN/STEP_A/tmp2[1] ), 
        .A(\MAIN/ENGIN/STEP_A/n3548 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U214  ( .ZN(\MAIN/ENGIN/STEP_A/n3577 ), .A(
        \MAIN/ENGIN/STEP_A/cst[1] ), .B(\MAIN/ENGIN/STEP_A/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/U221  ( .ZN(\MAIN/ENGIN/STEP_A/n3544 ), .A(
        \MAIN/ENGIN/STEP_A/cst[2] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_A/U233  ( .ZN(\MAIN/ENGIN/STEP_A/n3558 ), 
        .A(\MAIN/ENGIN/STEP_A/sw_stage ), .B(\MAIN/sw_end ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_A/U246  ( .ZN(\MAIN/ENGIN/STEP_A/n3551 ), .A(
        \MAIN/ENGIN/STEP_A/n3589 ), .B(\MAIN/ENGIN/STEP_A/n3563 ) );
    snl_aoi023x0 \MAIN/ENGIN/STEP_A/U228  ( .ZN(\MAIN/ENGIN/STEP_A/n3575 ), 
        .A(\MAIN/ENGIN/cf_start ), .B(\MAIN/ENGIN/STEP_A/n3568 ), .C(
        \MAIN/ENGIN/STEP_A/n3569 ), .D(\MAIN/ENGIN/STEP_A/d3_stage ), .E(
        \MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U191  ( .ZN(\MAIN/ENGIN/STEP_B/tmp2[0] ), 
        .A(\MAIN/ENGIN/STEP_B/n3498 ), .B(\MAIN/ENGIN/STEP_B/n3499 ) );
    snl_oai113x0 \MAIN/ENGIN/STEP_B/U198  ( .ZN(\MAIN/ENGIN/b_swctl_st ), .A(
        \MAIN/ENGIN/STEP_B/n3496 ), .B(\MAIN/exe_end ), .C(
        \MAIN/ENGIN/STEP_B/n3515 ), .D(\MAIN/ENGIN/STEP_B/n3516 ), .E(
        \MAIN/ENGIN/STEP_B/n3517 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_B/U204  ( .ZN(
        \MAIN/ENGIN/STEP_B/decode_stage272 ), .A(\MAIN/ENGIN/STEP_B/n3519 ), 
        .B(\MAIN/ENGIN/STEP_B/tmp2[2] ), .C(\MAIN/ENGIN/STEP_B/n3500 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_B/U223  ( .ZN(\MAIN/ENGIN/STEP_B/n3532 ), 
        .A(\MAIN/ENGIN/STEP_B/cst[0] ), .B(\MAIN/ENGIN/STEP_B/n3523 ), .C(
        \MAIN/ENGIN/STEP_B/n3529 ) );
    snl_aoi222x0 \MAIN/ENGIN/STEP_B/U238  ( .ZN(\MAIN/ENGIN/STEP_B/n3517 ), 
        .A(\MAIN/ENGIN/B_INIT_STAGE ), .B(\MAIN/ENGIN/STEP_B/n3530 ), .C(
        \MAIN/ENGIN/STEP_B/n3529 ), .D(\MAIN/ENGIN/STEP_B/n3528 ), .E(
        \MAIN/ENGIN/STEP_B/n3539 ), .F(\MAIN/ENGIN/STEP_B/n3523 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_B/U256  ( .ZN(\MAIN/ENGIN/STEP_B/n3537 ), 
        .A(\MAIN/ENGIN/STEP_B/n3509 ), .B(\MAIN/ENGIN/STEP_B/n3534 ), .C(
        \MAIN/ENGIN/STEP_B/n3527 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U196  ( .ZN(\MAIN/ENGIN/b_decctl_st ), .A(
        \MAIN/ENGIN/STEP_B/n3513 ), .B(\MAIN/ENGIN/STEP_B/n3514 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U211  ( .ZN(\MAIN/ENGIN/STEP_B/n3515 ), 
        .A(\MAIN/ENGIN/STEP_B/cst[1] ), .B(\MAIN/ENGIN/STEP_B/cst[0] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U216  ( .ZN(\MAIN/ENGIN/STEP_B/n3531 ), 
        .A(\MAIN/ENGIN/STEP_B/n3529 ), .B(\MAIN/ENGIN/STEP_B/n3521 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_B/U231  ( .ZN(\MAIN/ENGIN/STEP_B/n3526 ), .A(
        \MAIN/ENGIN/STEP_B/cst[2] ), .B(\MAIN/ENGIN/STEP_B/cst[3] ), .C(
        \MAIN/ENGIN/STEP_B/n3520 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U244  ( .ZN(\MAIN/ENGIN/STEP_B/cf_st2_rst ), 
        .A(\MAIN/ENGIN/STEP_B/n3533 ) );
    snl_aoi122x0 \MAIN/ENGIN/STEP_B/U236  ( .ZN(\MAIN/ENGIN/STEP_B/n3498 ), 
        .A(pk_pexe01_h), .B(\MAIN/ENGIN/STEP_B/n3537 ), .C(
        \MAIN/ENGIN/STEP_B/n3508 ), .D(\MAIN/ENGIN/STEP_B/n3538 ), .E(
        \MAIN/ENGIN/STEP_B/n3507 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U243  ( .ZN(step2_cf), .A(
        \MAIN/ENGIN/STEP_B/n3533 ), .B(pgperrh) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U258  ( .ZN(\MAIN/ENGIN/STEP_B/n3519 ), .A(
        \MAIN/ENGIN/STEP_B/tmp2[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U218  ( .ZN(\MAIN/ENGIN/STEP_B/n3512 ), .A(
        pk_pexe01_h) );
    snl_ao1b1b3x0 \MAIN/ENGIN/STEP_B/U251  ( .Z(\MAIN/ENGIN/STEP_B/n3505 ), 
        .A(\MAIN/ENGIN/STEP_B/n3540 ), .B(\MAIN/ENGIN/a_decctl_st ), .C(
        \MAIN/excep_valid ), .D(\MAIN/ENGIN/STEP_B/n3520 ), .E(
        \MAIN/ENGIN/STEP_B/n3542 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U190  ( .ZN(\MAIN/ENGIN/b_d2_stage ), .A(
        \MAIN/ENGIN/STEP_B/n3496 ), .B(\MAIN/ENGIN/STEP_B/n3497 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_B/U197  ( .ZN(\MAIN/ENGIN/b_exectl_st ), .A(
        \MAIN/ENGIN/STEP_B/n3508 ), .B(\MAIN/ENGIN/STEP_B/n3496 ), .C(
        \MAIN/ENGIN/STEP_B/n3506 ) );
    snl_ao112x1 \MAIN/ENGIN/STEP_B/U203  ( .Z(\MAIN/ENGIN/c_dec_start ), .A(
        \MAIN/ENGIN/STEP_B/n3520 ), .B(\MAIN/ENGIN/STEP_B/n3521 ), .C(
        \MAIN/ENGIN/STEP_B/n3506 ), .D(\MAIN/ENGIN/STEP_B/cst[2] ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_B/U224  ( .ZN(\MAIN/ENGIN/STEP_B/n3533 ), 
        .A(\MAIN/ENGIN/b_cf_stage ), .B(\MAIN/ENGIN/STEP_B/n3508 ), .C(
        pgiaendp) );
    snl_aoi112x0 \MAIN/ENGIN/STEP_B/U199  ( .ZN(
        \MAIN/ENGIN/STEP_B/dec_st2_rst ), .A(\MAIN/ENGIN/STEP_B/n3508 ), .B(
        \MAIN/ENGIN/STEP_B/n3518 ), .C(\MAIN/ENGIN/STEP_B/n3515 ), .D(
        \MAIN/ENGIN/STEP_B/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U202  ( .ZN(ph_dec_bh), .A(
        \MAIN/ENGIN/b_dec_stage ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U210  ( .ZN(\MAIN/ENGIN/STEP_B/n3520 ), .A(
        \MAIN/ENGIN/STEP_B/cst[1] ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U242  ( .ZN(\MAIN/ENGIN/b_step_end ), .A(
        \MAIN/ENGIN/STEP_B/n3510 ) );
    snl_ao022x1 \MAIN/ENGIN/STEP_B/U259  ( .Z(\MAIN/ENGIN/STEP_B/n3541 ), .A(
        \MAIN/exe_end ), .B(\MAIN/ENGIN/STEP_B/cst[2] ), .C(
        \MAIN/ENGIN/STEP_B/n3535 ), .D(\MAIN/ENGIN/STEP_B/n3496 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_B/cst_reg[0]  ( .Q(\MAIN/ENGIN/STEP_B/cst[0] 
        ), .D(\MAIN/ENGIN/STEP_B/tmp2[0] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U237  ( .ZN(\MAIN/ENGIN/STEP_B/n3516 ), .A(
        \MAIN/ENGIN/STEP_B/n3526 ), .B(\MAIN/ENGIN/STEP_B/n3502 ) );
    snl_and34x0 \MAIN/ENGIN/STEP_B/U205  ( .Z(\MAIN/ENGIN/STEP_B/n3522 ), .A(
        \MAIN/ENGIN/STEP_B/cst[1] ), .B(\MAIN/ENGIN/STEP_B/cst[0] ), .C(
        \MAIN/ENGIN/STEP_B/n3523 ), .D(\MAIN/POL_STH ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U219  ( .ZN(\MAIN/ENGIN/STEP_B/n3508 ), .A(
        \MAIN/ENGIN/STEP_B/n3512 ), .B(\MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U225  ( .ZN(\MAIN/ENGIN/STEP_B/n3534 ), 
        .A(\MAIN/ENGIN/STEP_B/cst[2] ), .B(\MAIN/ENGIN/STEP_B/n3520 ) );
    snl_aoi012x1 \MAIN/ENGIN/STEP_B/U250  ( .ZN(\MAIN/ENGIN/STEP_B/n3542 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/a_decctl_st ), .C(
        \MAIN/ENGIN/STEP_B/n3525 ) );
    snl_ao01b2x0 \MAIN/ENGIN/STEP_B/U222  ( .Z(\MAIN/ENGIN/STEP_B/n3507 ), .A(
        \MAIN/ENGIN/STEP_B/n3530 ), .B(\MAIN/ENGIN/STEP_B/n3531 ), .C(
        \MAIN/ENGIN/status_wr2 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U239  ( .ZN(\MAIN/ENGIN/B_INIT_STAGE ), .A(
        \MAIN/ENGIN/STEP_B/n3531 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U257  ( .ZN(\MAIN/ENGIN/STEP_B/n3536 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/STEP_B/n3509 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U217  ( .ZN(\MAIN/ENGIN/STEP_B/n3523 ), .A(
        \MAIN/ENGIN/STEP_B/cst[3] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U230  ( .ZN(\MAIN/ENGIN/STEP_B/n3506 ), .A(
        \MAIN/ENGIN/STEP_B/n3518 ), .B(\MAIN/ENGIN/STEP_B/n3515 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U245  ( .ZN(\MAIN/ENGIN/STEP_B/n3540 ), .A(
        \MAIN/ENGIN/STEP_B/n3508 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_B/cst_reg[2]  ( .Q(\MAIN/ENGIN/STEP_B/cst[2] 
        ), .D(\MAIN/ENGIN/STEP_B/tmp2[2] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_B/exec_stage_reg  ( .Q(\MAIN/b_exec_stage ), 
        .D(\MAIN/ENGIN/STEP_B/exec_stage278 ), .RN(\MAIN/ENGIN/n3591 ), .CP(
        SCLK) );
    snl_and34x0 \MAIN/ENGIN/STEP_B/U192  ( .Z(\MAIN/ENGIN/STEP_B/n3500 ), .A(
        \MAIN/ENGIN/STEP_B/n3502 ), .B(\MAIN/ENGIN/STEP_B/n3503 ), .C(step2_cf
        ), .D(\MAIN/ENGIN/STEP_B/n3501 ) );
    snl_aoi013x0 \MAIN/ENGIN/STEP_B/U207  ( .ZN(\MAIN/ENGIN/STEP_B/n3513 ), 
        .A(\MAIN/ENGIN/STEP_B/n3508 ), .B(\MAIN/ENGIN/STEP_B/n3525 ), .C(
        \MAIN/ENGIN/STEP_B/n3526 ), .D(step2_cf) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U220  ( .ZN(\MAIN/ENGIN/STEP_B/n3509 ), .A(
        \MAIN/ENGIN/a_decctl_st ) );
    snl_oai233x0 \MAIN/ENGIN/STEP_B/U255  ( .ZN(\MAIN/ENGIN/STEP_B/n3538 ), 
        .A(\MAIN/ENGIN/STEP_B/n3523 ), .B(\MAIN/ENGIN/B_PED4_BR ), .C(
        \MAIN/ENGIN/STEP_B/n3525 ), .D(\MAIN/ENGIN/STEP_B/n3514 ), .E(
        \MAIN/ENGIN/STEP_B/cst[2] ), .F(\MAIN/ENGIN/STEP_B/n3520 ), .G(
        \MAIN/ENGIN/STEP_B/n3524 ), .H(\MAIN/ENGIN/STEP_B/n3532 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_B/cst_reg[3]  ( .Q(\MAIN/ENGIN/STEP_B/cst[3] 
        ), .D(\MAIN/ENGIN/STEP_B/nst[3] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_B/U193  ( .ZN(\MAIN/ENGIN/STEP_B/n3504 ), 
        .A(\MAIN/ENGIN/STEP_B/cst[2] ), .B(\MAIN/ENGIN/STEP_B/n3505 ), .C(
        \MAIN/ENGIN/STEP_B/n3506 ), .D(\MAIN/ENGIN/STEP_B/n3507 ) );
    snl_ao023x1 \MAIN/ENGIN/STEP_B/U194  ( .Z(\MAIN/ENGIN/STEP_B/nst[3] ), .A(
        \MAIN/ENGIN/STEP_B/n3508 ), .B(\MAIN/ENGIN/STEP_B/n3497 ), .C(
        \MAIN/ENGIN/STEP_B/cst[3] ), .D(\MAIN/ENGIN/STEP_B/cf_st2_rst ), .E(
        pgperrh) );
    snl_oai022x1 \MAIN/ENGIN/STEP_B/U195  ( .ZN(\MAIN/ENGIN/b_cfctl_st ), .A(
        \MAIN/ENGIN/STEP_B/n3509 ), .B(\MAIN/ENGIN/STEP_B/n3510 ), .C(
        \MAIN/ENGIN/STEP_B/n3511 ), .D(\MAIN/ENGIN/STEP_B/n3512 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U212  ( .ZN(\MAIN/ENGIN/STEP_B/n3518 ), .A(
        \MAIN/dec_end ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_B/U215  ( .ZN(\MAIN/ENGIN/STEP_B/n3530 ), 
        .A(\MAIN/ENGIN/STEP_B/n3509 ), .B(\MAIN/ENGIN/STEP_B/n3512 ), .C(
        \MAIN/POL_STH ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U229  ( .ZN(\MAIN/ENGIN/STEP_B/n3514 ), .A(
        \MAIN/ENGIN/b_dec_start ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_B/decode_stage_reg  ( .Q(
        \MAIN/ENGIN/b_dec_stage ), .D(\MAIN/ENGIN/STEP_B/decode_stage272 ), 
        .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK) );
    snl_nor03x0 \MAIN/ENGIN/STEP_B/U247  ( .ZN(\MAIN/ENGIN/STEP_B/n3502 ), .A(
        \MAIN/ENGIN/STEP_B/n3520 ), .B(pol_status), .C(
        \MAIN/ENGIN/STEP_B/n3496 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U232  ( .ZN(\MAIN/ENGIN/STEP_B/n3497 ), 
        .A(\MAIN/ENGIN/STEP_B/cst[1] ), .B(\MAIN/ENGIN/STEP_B/n3525 ) );
    snl_aoi123x0 \MAIN/ENGIN/STEP_B/U235  ( .ZN(\MAIN/ENGIN/STEP_B/n3499 ), 
        .A(\MAIN/ENGIN/STEP_B/cst[2] ), .B(\MAIN/ENGIN/STEP_B/cst[1] ), .C(
        pol_status), .D(\MAIN/ENGIN/STEP_B/sw_stage ), .E(
        \MAIN/ENGIN/STEP_B/n3536 ), .F(\MAIN/ENGIN/STEP_B/n3503 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U240  ( .ZN(\MAIN/ENGIN/b_cf_stage ), .A(
        \MAIN/ENGIN/STEP_B/n3532 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_B/U200  ( .ZN(
        \MAIN/ENGIN/STEP_B/exec_stage278 ), .A(\MAIN/ENGIN/STEP_B/n3519 ), .B(
        \MAIN/ENGIN/STEP_B/n3504 ), .C(\MAIN/ENGIN/STEP_B/n3500 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U209  ( .ZN(\MAIN/ENGIN/STEP_B/n3525 ), .A(
        \MAIN/ENGIN/STEP_B/cst[0] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U227  ( .ZN(\MAIN/ENGIN/STEP_B/d3_stage ), 
        .A(\MAIN/ENGIN/STEP_B/n3534 ), .B(\MAIN/ENGIN/STEP_B/cst[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U249  ( .ZN(\MAIN/ENGIN/STEP_B/n3521 ), .A(
        \MAIN/ENGIN/STEP_B/n3528 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U252  ( .ZN(\MAIN/ENGIN/STEP_B/tmp2[2] ), 
        .A(\MAIN/ENGIN/STEP_B/n3504 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_B/cst_reg[1]  ( .Q(\MAIN/ENGIN/STEP_B/cst[1] 
        ), .D(\MAIN/ENGIN/STEP_B/tmp2[1] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_invx05 \MAIN/ENGIN/STEP_B/U201  ( .ZN(ph_exe_bh), .A(
        \MAIN/b_exec_stage ) );
    snl_aoi0b12x0 \MAIN/ENGIN/STEP_B/U208  ( .ZN(\MAIN/ENGIN/STEP_B/n3511 ), 
        .A(\MAIN/ENGIN/STEP_B/d3_stage ), .B(\MAIN/ENGIN/a_decctl_st ), .C(
        \MAIN/ENGIN/STEP_B/n3527 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U213  ( .ZN(\MAIN/ENGIN/STEP_B/n3528 ), 
        .A(\MAIN/ENGIN/STEP_B/n3523 ), .B(\MAIN/ENGIN/STEP_B/n3525 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U234  ( .ZN(\MAIN/ENGIN/STEP_B/n3535 ), .A(
        \MAIN/dec_end ), .B(\MAIN/ENGIN/STEP_B/n3508 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U241  ( .ZN(\MAIN/ENGIN/status_wr2 ), .A(
        \MAIN/ENGIN/STEP_B/n3523 ), .B(\MAIN/ENGIN/STEP_B/n3520 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U226  ( .ZN(\MAIN/ENGIN/STEP_B/sw_stage ), 
        .A(\MAIN/ENGIN/STEP_B/n3534 ), .B(\MAIN/ENGIN/STEP_B/n3525 ) );
    snl_and23x0 \MAIN/ENGIN/STEP_B/U206  ( .Z(\MAIN/ENGIN/STEP_B/n3524 ), .A(
        \MAIN/ENGIN/b_dec_start ), .B(pgperrh), .C(pgiaendp) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U248  ( .ZN(\MAIN/ENGIN/STEP_B/n3539 ), .A(
        \MAIN/ENGIN/STEP_B/n3534 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_B/U253  ( .ZN(\MAIN/ENGIN/STEP_B/n3501 ), 
        .A(\MAIN/ENGIN/STEP_B/n3522 ), .B(\MAIN/ENGIN/STEP_B/n3526 ), .C(
        \MAIN/ENGIN/STEP_B/n3508 ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U254  ( .ZN(\MAIN/ENGIN/STEP_B/tmp2[1] ), 
        .A(\MAIN/ENGIN/STEP_B/n3500 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U214  ( .ZN(\MAIN/ENGIN/STEP_B/n3529 ), .A(
        \MAIN/ENGIN/STEP_B/cst[1] ), .B(\MAIN/ENGIN/STEP_B/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/U221  ( .ZN(\MAIN/ENGIN/STEP_B/n3496 ), .A(
        \MAIN/ENGIN/STEP_B/cst[2] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_B/U233  ( .ZN(\MAIN/ENGIN/STEP_B/n3510 ), 
        .A(\MAIN/ENGIN/STEP_B/sw_stage ), .B(\MAIN/sw_end ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_B/U246  ( .ZN(\MAIN/ENGIN/STEP_B/n3503 ), .A(
        \MAIN/ENGIN/STEP_B/n3541 ), .B(\MAIN/ENGIN/STEP_B/n3515 ) );
    snl_aoi023x0 \MAIN/ENGIN/STEP_B/U228  ( .ZN(\MAIN/ENGIN/STEP_B/n3527 ), 
        .A(\MAIN/ENGIN/a_decctl_st ), .B(\MAIN/ENGIN/STEP_B/n3520 ), .C(
        \MAIN/ENGIN/STEP_B/n3521 ), .D(\MAIN/ENGIN/STEP_B/d3_stage ), .E(
        \MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U191  ( .ZN(\MAIN/ENGIN/STEP_C/tmp2[0] ), 
        .A(\MAIN/ENGIN/STEP_C/n3450 ), .B(\MAIN/ENGIN/STEP_C/n3451 ) );
    snl_oai113x0 \MAIN/ENGIN/STEP_C/U198  ( .ZN(\MAIN/ENGIN/c_swctl_st ), .A(
        \MAIN/ENGIN/STEP_C/n3448 ), .B(\MAIN/exe_end ), .C(
        \MAIN/ENGIN/STEP_C/n3467 ), .D(\MAIN/ENGIN/STEP_C/n3468 ), .E(
        \MAIN/ENGIN/STEP_C/n3469 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_C/U204  ( .ZN(
        \MAIN/ENGIN/STEP_C/decode_stage272 ), .A(\MAIN/ENGIN/STEP_C/n3471 ), 
        .B(\MAIN/ENGIN/STEP_C/tmp2[2] ), .C(\MAIN/ENGIN/STEP_C/n3452 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_C/U223  ( .ZN(\MAIN/ENGIN/STEP_C/n3484 ), 
        .A(\MAIN/ENGIN/STEP_C/cst[0] ), .B(\MAIN/ENGIN/STEP_C/n3475 ), .C(
        \MAIN/ENGIN/STEP_C/n3481 ) );
    snl_aoi222x0 \MAIN/ENGIN/STEP_C/U238  ( .ZN(\MAIN/ENGIN/STEP_C/n3469 ), 
        .A(\MAIN/ENGIN/C_INIT_STAGE ), .B(\MAIN/ENGIN/STEP_C/n3482 ), .C(
        \MAIN/ENGIN/STEP_C/n3481 ), .D(\MAIN/ENGIN/STEP_C/n3480 ), .E(
        \MAIN/ENGIN/STEP_C/n3491 ), .F(\MAIN/ENGIN/STEP_C/n3475 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_C/U256  ( .ZN(\MAIN/ENGIN/STEP_C/n3489 ), 
        .A(\MAIN/ENGIN/STEP_C/n3461 ), .B(\MAIN/ENGIN/STEP_C/n3486 ), .C(
        \MAIN/ENGIN/STEP_C/n3479 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U196  ( .ZN(\MAIN/ENGIN/c_decctl_st ), .A(
        \MAIN/ENGIN/STEP_C/n3465 ), .B(\MAIN/ENGIN/STEP_C/n3466 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U211  ( .ZN(\MAIN/ENGIN/STEP_C/n3467 ), 
        .A(\MAIN/ENGIN/STEP_C/cst[1] ), .B(\MAIN/ENGIN/STEP_C/cst[0] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U216  ( .ZN(\MAIN/ENGIN/STEP_C/n3483 ), 
        .A(\MAIN/ENGIN/STEP_C/n3481 ), .B(\MAIN/ENGIN/STEP_C/n3473 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_C/U231  ( .ZN(\MAIN/ENGIN/STEP_C/n3478 ), .A(
        \MAIN/ENGIN/STEP_C/cst[2] ), .B(\MAIN/ENGIN/STEP_C/cst[3] ), .C(
        \MAIN/ENGIN/STEP_C/n3472 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U244  ( .ZN(\MAIN/ENGIN/STEP_C/cf_st2_rst ), 
        .A(\MAIN/ENGIN/STEP_C/n3485 ) );
    snl_aoi122x0 \MAIN/ENGIN/STEP_C/U236  ( .ZN(\MAIN/ENGIN/STEP_C/n3450 ), 
        .A(pk_pexe01_h), .B(\MAIN/ENGIN/STEP_C/n3489 ), .C(
        \MAIN/ENGIN/STEP_C/n3460 ), .D(\MAIN/ENGIN/STEP_C/n3490 ), .E(
        \MAIN/ENGIN/STEP_C/n3459 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U243  ( .ZN(step3_cf), .A(
        \MAIN/ENGIN/STEP_C/n3485 ), .B(pgperrh) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U258  ( .ZN(\MAIN/ENGIN/STEP_C/n3471 ), .A(
        \MAIN/ENGIN/STEP_C/tmp2[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U218  ( .ZN(\MAIN/ENGIN/STEP_C/n3464 ), .A(
        pk_pexe01_h) );
    snl_ao1b1b3x0 \MAIN/ENGIN/STEP_C/U251  ( .Z(\MAIN/ENGIN/STEP_C/n3457 ), 
        .A(\MAIN/ENGIN/STEP_C/n3492 ), .B(\MAIN/ENGIN/b_decctl_st ), .C(
        \MAIN/excep_valid ), .D(\MAIN/ENGIN/STEP_C/n3472 ), .E(
        \MAIN/ENGIN/STEP_C/n3494 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U190  ( .ZN(\MAIN/ENGIN/c_d2_stage ), .A(
        \MAIN/ENGIN/STEP_C/n3448 ), .B(\MAIN/ENGIN/STEP_C/n3449 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_C/U197  ( .ZN(\MAIN/ENGIN/c_exectl_st ), .A(
        \MAIN/ENGIN/STEP_C/n3460 ), .B(\MAIN/ENGIN/STEP_C/n3448 ), .C(
        \MAIN/ENGIN/STEP_C/n3458 ) );
    snl_ao112x1 \MAIN/ENGIN/STEP_C/U203  ( .Z(\MAIN/ENGIN/d_dec_start ), .A(
        \MAIN/ENGIN/STEP_C/n3472 ), .B(\MAIN/ENGIN/STEP_C/n3473 ), .C(
        \MAIN/ENGIN/STEP_C/n3458 ), .D(\MAIN/ENGIN/STEP_C/cst[2] ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_C/U224  ( .ZN(\MAIN/ENGIN/STEP_C/n3485 ), 
        .A(\MAIN/ENGIN/c_cf_stage ), .B(\MAIN/ENGIN/STEP_C/n3460 ), .C(
        pgiaendp) );
    snl_aoi112x0 \MAIN/ENGIN/STEP_C/U199  ( .ZN(
        \MAIN/ENGIN/STEP_C/dec_st2_rst ), .A(\MAIN/ENGIN/STEP_C/n3460 ), .B(
        \MAIN/ENGIN/STEP_C/n3470 ), .C(\MAIN/ENGIN/STEP_C/n3467 ), .D(
        \MAIN/ENGIN/STEP_C/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U202  ( .ZN(ph_dec_ch), .A(
        \MAIN/ENGIN/c_dec_stage ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U210  ( .ZN(\MAIN/ENGIN/STEP_C/n3472 ), .A(
        \MAIN/ENGIN/STEP_C/cst[1] ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U242  ( .ZN(\MAIN/ENGIN/c_step_end ), .A(
        \MAIN/ENGIN/STEP_C/n3462 ) );
    snl_ao022x1 \MAIN/ENGIN/STEP_C/U259  ( .Z(\MAIN/ENGIN/STEP_C/n3493 ), .A(
        \MAIN/exe_end ), .B(\MAIN/ENGIN/STEP_C/cst[2] ), .C(
        \MAIN/ENGIN/STEP_C/n3487 ), .D(\MAIN/ENGIN/STEP_C/n3448 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_C/cst_reg[0]  ( .Q(\MAIN/ENGIN/STEP_C/cst[0] 
        ), .D(\MAIN/ENGIN/STEP_C/tmp2[0] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U237  ( .ZN(\MAIN/ENGIN/STEP_C/n3468 ), .A(
        \MAIN/ENGIN/STEP_C/n3478 ), .B(\MAIN/ENGIN/STEP_C/n3454 ) );
    snl_and34x0 \MAIN/ENGIN/STEP_C/U205  ( .Z(\MAIN/ENGIN/STEP_C/n3474 ), .A(
        \MAIN/ENGIN/STEP_C/cst[1] ), .B(\MAIN/ENGIN/STEP_C/cst[0] ), .C(
        \MAIN/ENGIN/STEP_C/n3475 ), .D(\MAIN/POL_STH ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U219  ( .ZN(\MAIN/ENGIN/STEP_C/n3460 ), .A(
        \MAIN/ENGIN/STEP_C/n3464 ), .B(\MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U225  ( .ZN(\MAIN/ENGIN/STEP_C/n3486 ), 
        .A(\MAIN/ENGIN/STEP_C/cst[2] ), .B(\MAIN/ENGIN/STEP_C/n3472 ) );
    snl_aoi012x1 \MAIN/ENGIN/STEP_C/U250  ( .ZN(\MAIN/ENGIN/STEP_C/n3494 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/b_decctl_st ), .C(
        \MAIN/ENGIN/STEP_C/n3477 ) );
    snl_ao01b2x0 \MAIN/ENGIN/STEP_C/U222  ( .Z(\MAIN/ENGIN/STEP_C/n3459 ), .A(
        \MAIN/ENGIN/STEP_C/n3482 ), .B(\MAIN/ENGIN/STEP_C/n3483 ), .C(
        \MAIN/ENGIN/status_wr3 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U239  ( .ZN(\MAIN/ENGIN/C_INIT_STAGE ), .A(
        \MAIN/ENGIN/STEP_C/n3483 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U257  ( .ZN(\MAIN/ENGIN/STEP_C/n3488 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/STEP_C/n3461 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U217  ( .ZN(\MAIN/ENGIN/STEP_C/n3475 ), .A(
        \MAIN/ENGIN/STEP_C/cst[3] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U230  ( .ZN(\MAIN/ENGIN/STEP_C/n3458 ), .A(
        \MAIN/ENGIN/STEP_C/n3470 ), .B(\MAIN/ENGIN/STEP_C/n3467 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U245  ( .ZN(\MAIN/ENGIN/STEP_C/n3492 ), .A(
        \MAIN/ENGIN/STEP_C/n3460 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_C/cst_reg[2]  ( .Q(\MAIN/ENGIN/STEP_C/cst[2] 
        ), .D(\MAIN/ENGIN/STEP_C/tmp2[2] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_C/exec_stage_reg  ( .Q(\MAIN/c_exec_stage ), 
        .D(\MAIN/ENGIN/STEP_C/exec_stage278 ), .RN(\MAIN/ENGIN/n3591 ), .CP(
        SCLK) );
    snl_and34x0 \MAIN/ENGIN/STEP_C/U192  ( .Z(\MAIN/ENGIN/STEP_C/n3452 ), .A(
        \MAIN/ENGIN/STEP_C/n3454 ), .B(\MAIN/ENGIN/STEP_C/n3455 ), .C(step3_cf
        ), .D(\MAIN/ENGIN/STEP_C/n3453 ) );
    snl_aoi013x0 \MAIN/ENGIN/STEP_C/U207  ( .ZN(\MAIN/ENGIN/STEP_C/n3465 ), 
        .A(\MAIN/ENGIN/STEP_C/n3460 ), .B(\MAIN/ENGIN/STEP_C/n3477 ), .C(
        \MAIN/ENGIN/STEP_C/n3478 ), .D(step3_cf) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U220  ( .ZN(\MAIN/ENGIN/STEP_C/n3461 ), .A(
        \MAIN/ENGIN/b_decctl_st ) );
    snl_oai233x0 \MAIN/ENGIN/STEP_C/U255  ( .ZN(\MAIN/ENGIN/STEP_C/n3490 ), 
        .A(\MAIN/ENGIN/STEP_C/n3475 ), .B(\MAIN/ENGIN/C_PED4_BR ), .C(
        \MAIN/ENGIN/STEP_C/n3477 ), .D(\MAIN/ENGIN/STEP_C/n3466 ), .E(
        \MAIN/ENGIN/STEP_C/cst[2] ), .F(\MAIN/ENGIN/STEP_C/n3472 ), .G(
        \MAIN/ENGIN/STEP_C/n3476 ), .H(\MAIN/ENGIN/STEP_C/n3484 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_C/cst_reg[3]  ( .Q(\MAIN/ENGIN/STEP_C/cst[3] 
        ), .D(\MAIN/ENGIN/STEP_C/nst[3] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_C/U193  ( .ZN(\MAIN/ENGIN/STEP_C/n3456 ), 
        .A(\MAIN/ENGIN/STEP_C/cst[2] ), .B(\MAIN/ENGIN/STEP_C/n3457 ), .C(
        \MAIN/ENGIN/STEP_C/n3458 ), .D(\MAIN/ENGIN/STEP_C/n3459 ) );
    snl_ao023x1 \MAIN/ENGIN/STEP_C/U194  ( .Z(\MAIN/ENGIN/STEP_C/nst[3] ), .A(
        \MAIN/ENGIN/STEP_C/n3460 ), .B(\MAIN/ENGIN/STEP_C/n3449 ), .C(
        \MAIN/ENGIN/STEP_C/cst[3] ), .D(\MAIN/ENGIN/STEP_C/cf_st2_rst ), .E(
        pgperrh) );
    snl_oai022x1 \MAIN/ENGIN/STEP_C/U195  ( .ZN(\MAIN/ENGIN/c_cfctl_st ), .A(
        \MAIN/ENGIN/STEP_C/n3461 ), .B(\MAIN/ENGIN/STEP_C/n3462 ), .C(
        \MAIN/ENGIN/STEP_C/n3463 ), .D(\MAIN/ENGIN/STEP_C/n3464 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U212  ( .ZN(\MAIN/ENGIN/STEP_C/n3470 ), .A(
        \MAIN/dec_end ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_C/U215  ( .ZN(\MAIN/ENGIN/STEP_C/n3482 ), 
        .A(\MAIN/ENGIN/STEP_C/n3461 ), .B(\MAIN/ENGIN/STEP_C/n3464 ), .C(
        \MAIN/POL_STH ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U229  ( .ZN(\MAIN/ENGIN/STEP_C/n3466 ), .A(
        \MAIN/ENGIN/c_dec_start ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_C/decode_stage_reg  ( .Q(
        \MAIN/ENGIN/c_dec_stage ), .D(\MAIN/ENGIN/STEP_C/decode_stage272 ), 
        .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK) );
    snl_nor03x0 \MAIN/ENGIN/STEP_C/U247  ( .ZN(\MAIN/ENGIN/STEP_C/n3454 ), .A(
        \MAIN/ENGIN/STEP_C/n3472 ), .B(pol_status), .C(
        \MAIN/ENGIN/STEP_C/n3448 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U232  ( .ZN(\MAIN/ENGIN/STEP_C/n3449 ), 
        .A(\MAIN/ENGIN/STEP_C/cst[1] ), .B(\MAIN/ENGIN/STEP_C/n3477 ) );
    snl_aoi123x0 \MAIN/ENGIN/STEP_C/U235  ( .ZN(\MAIN/ENGIN/STEP_C/n3451 ), 
        .A(\MAIN/ENGIN/STEP_C/cst[2] ), .B(\MAIN/ENGIN/STEP_C/cst[1] ), .C(
        pol_status), .D(\MAIN/ENGIN/STEP_C/sw_stage ), .E(
        \MAIN/ENGIN/STEP_C/n3488 ), .F(\MAIN/ENGIN/STEP_C/n3455 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U240  ( .ZN(\MAIN/ENGIN/c_cf_stage ), .A(
        \MAIN/ENGIN/STEP_C/n3484 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_C/U200  ( .ZN(
        \MAIN/ENGIN/STEP_C/exec_stage278 ), .A(\MAIN/ENGIN/STEP_C/n3471 ), .B(
        \MAIN/ENGIN/STEP_C/n3456 ), .C(\MAIN/ENGIN/STEP_C/n3452 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U209  ( .ZN(\MAIN/ENGIN/STEP_C/n3477 ), .A(
        \MAIN/ENGIN/STEP_C/cst[0] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U227  ( .ZN(\MAIN/ENGIN/STEP_C/d3_stage ), 
        .A(\MAIN/ENGIN/STEP_C/n3486 ), .B(\MAIN/ENGIN/STEP_C/cst[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U249  ( .ZN(\MAIN/ENGIN/STEP_C/n3473 ), .A(
        \MAIN/ENGIN/STEP_C/n3480 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U252  ( .ZN(\MAIN/ENGIN/STEP_C/tmp2[2] ), 
        .A(\MAIN/ENGIN/STEP_C/n3456 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_C/cst_reg[1]  ( .Q(\MAIN/ENGIN/STEP_C/cst[1] 
        ), .D(\MAIN/ENGIN/STEP_C/tmp2[1] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_invx05 \MAIN/ENGIN/STEP_C/U201  ( .ZN(ph_exe_ch), .A(
        \MAIN/c_exec_stage ) );
    snl_aoi0b12x0 \MAIN/ENGIN/STEP_C/U208  ( .ZN(\MAIN/ENGIN/STEP_C/n3463 ), 
        .A(\MAIN/ENGIN/STEP_C/d3_stage ), .B(\MAIN/ENGIN/b_decctl_st ), .C(
        \MAIN/ENGIN/STEP_C/n3479 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U213  ( .ZN(\MAIN/ENGIN/STEP_C/n3480 ), 
        .A(\MAIN/ENGIN/STEP_C/n3475 ), .B(\MAIN/ENGIN/STEP_C/n3477 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U234  ( .ZN(\MAIN/ENGIN/STEP_C/n3487 ), .A(
        \MAIN/dec_end ), .B(\MAIN/ENGIN/STEP_C/n3460 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U241  ( .ZN(\MAIN/ENGIN/status_wr3 ), .A(
        \MAIN/ENGIN/STEP_C/n3475 ), .B(\MAIN/ENGIN/STEP_C/n3472 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U226  ( .ZN(\MAIN/ENGIN/STEP_C/sw_stage ), 
        .A(\MAIN/ENGIN/STEP_C/n3486 ), .B(\MAIN/ENGIN/STEP_C/n3477 ) );
    snl_and23x0 \MAIN/ENGIN/STEP_C/U206  ( .Z(\MAIN/ENGIN/STEP_C/n3476 ), .A(
        \MAIN/ENGIN/c_dec_start ), .B(pgperrh), .C(pgiaendp) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U248  ( .ZN(\MAIN/ENGIN/STEP_C/n3491 ), .A(
        \MAIN/ENGIN/STEP_C/n3486 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_C/U253  ( .ZN(\MAIN/ENGIN/STEP_C/n3453 ), 
        .A(\MAIN/ENGIN/STEP_C/n3474 ), .B(\MAIN/ENGIN/STEP_C/n3478 ), .C(
        \MAIN/ENGIN/STEP_C/n3460 ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U254  ( .ZN(\MAIN/ENGIN/STEP_C/tmp2[1] ), 
        .A(\MAIN/ENGIN/STEP_C/n3452 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U214  ( .ZN(\MAIN/ENGIN/STEP_C/n3481 ), .A(
        \MAIN/ENGIN/STEP_C/cst[1] ), .B(\MAIN/ENGIN/STEP_C/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/U221  ( .ZN(\MAIN/ENGIN/STEP_C/n3448 ), .A(
        \MAIN/ENGIN/STEP_C/cst[2] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_C/U233  ( .ZN(\MAIN/ENGIN/STEP_C/n3462 ), 
        .A(\MAIN/ENGIN/STEP_C/sw_stage ), .B(\MAIN/sw_end ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_C/U246  ( .ZN(\MAIN/ENGIN/STEP_C/n3455 ), .A(
        \MAIN/ENGIN/STEP_C/n3493 ), .B(\MAIN/ENGIN/STEP_C/n3467 ) );
    snl_aoi023x0 \MAIN/ENGIN/STEP_C/U228  ( .ZN(\MAIN/ENGIN/STEP_C/n3479 ), 
        .A(\MAIN/ENGIN/b_decctl_st ), .B(\MAIN/ENGIN/STEP_C/n3472 ), .C(
        \MAIN/ENGIN/STEP_C/n3473 ), .D(\MAIN/ENGIN/STEP_C/d3_stage ), .E(
        \MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U191  ( .ZN(\MAIN/ENGIN/STEP_D/tmp2[0] ), 
        .A(\MAIN/ENGIN/STEP_D/n3402 ), .B(\MAIN/ENGIN/STEP_D/n3403 ) );
    snl_oai113x0 \MAIN/ENGIN/STEP_D/U198  ( .ZN(\MAIN/ENGIN/d_swctl_st ), .A(
        \MAIN/ENGIN/STEP_D/n3400 ), .B(\MAIN/exe_end ), .C(
        \MAIN/ENGIN/STEP_D/n3419 ), .D(\MAIN/ENGIN/STEP_D/n3420 ), .E(
        \MAIN/ENGIN/STEP_D/n3421 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_D/U204  ( .ZN(
        \MAIN/ENGIN/STEP_D/decode_stage272 ), .A(\MAIN/ENGIN/STEP_D/n3423 ), 
        .B(\MAIN/ENGIN/STEP_D/tmp2[2] ), .C(\MAIN/ENGIN/STEP_D/n3404 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_D/U223  ( .ZN(\MAIN/ENGIN/STEP_D/n3436 ), 
        .A(\MAIN/ENGIN/STEP_D/cst[0] ), .B(\MAIN/ENGIN/STEP_D/n3427 ), .C(
        \MAIN/ENGIN/STEP_D/n3433 ) );
    snl_aoi222x0 \MAIN/ENGIN/STEP_D/U238  ( .ZN(\MAIN/ENGIN/STEP_D/n3421 ), 
        .A(\MAIN/ENGIN/D_INIT_STAGE ), .B(\MAIN/ENGIN/STEP_D/n3434 ), .C(
        \MAIN/ENGIN/STEP_D/n3433 ), .D(\MAIN/ENGIN/STEP_D/n3432 ), .E(
        \MAIN/ENGIN/STEP_D/n3443 ), .F(\MAIN/ENGIN/STEP_D/n3427 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_D/U256  ( .ZN(\MAIN/ENGIN/STEP_D/n3441 ), 
        .A(\MAIN/ENGIN/STEP_D/n3413 ), .B(\MAIN/ENGIN/STEP_D/n3438 ), .C(
        \MAIN/ENGIN/STEP_D/n3431 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U196  ( .ZN(\MAIN/ENGIN/d_decctl_st ), .A(
        \MAIN/ENGIN/STEP_D/n3417 ), .B(\MAIN/ENGIN/STEP_D/n3418 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U211  ( .ZN(\MAIN/ENGIN/STEP_D/n3419 ), 
        .A(\MAIN/ENGIN/STEP_D/cst[1] ), .B(\MAIN/ENGIN/STEP_D/cst[0] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U216  ( .ZN(\MAIN/ENGIN/STEP_D/n3435 ), 
        .A(\MAIN/ENGIN/STEP_D/n3433 ), .B(\MAIN/ENGIN/STEP_D/n3425 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_D/U231  ( .ZN(\MAIN/ENGIN/STEP_D/n3430 ), .A(
        \MAIN/ENGIN/STEP_D/cst[2] ), .B(\MAIN/ENGIN/STEP_D/cst[3] ), .C(
        \MAIN/ENGIN/STEP_D/n3424 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U244  ( .ZN(\MAIN/ENGIN/STEP_D/cf_st2_rst ), 
        .A(\MAIN/ENGIN/STEP_D/n3437 ) );
    snl_aoi122x0 \MAIN/ENGIN/STEP_D/U236  ( .ZN(\MAIN/ENGIN/STEP_D/n3402 ), 
        .A(pk_pexe01_h), .B(\MAIN/ENGIN/STEP_D/n3441 ), .C(
        \MAIN/ENGIN/STEP_D/n3412 ), .D(\MAIN/ENGIN/STEP_D/n3442 ), .E(
        \MAIN/ENGIN/STEP_D/n3411 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U243  ( .ZN(step4_cf), .A(
        \MAIN/ENGIN/STEP_D/n3437 ), .B(pgperrh) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U258  ( .ZN(\MAIN/ENGIN/STEP_D/n3423 ), .A(
        \MAIN/ENGIN/STEP_D/tmp2[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U218  ( .ZN(\MAIN/ENGIN/STEP_D/n3416 ), .A(
        pk_pexe01_h) );
    snl_ao1b1b3x0 \MAIN/ENGIN/STEP_D/U251  ( .Z(\MAIN/ENGIN/STEP_D/n3409 ), 
        .A(\MAIN/ENGIN/STEP_D/n3444 ), .B(\MAIN/ENGIN/c_decctl_st ), .C(
        \MAIN/excep_valid ), .D(\MAIN/ENGIN/STEP_D/n3424 ), .E(
        \MAIN/ENGIN/STEP_D/n3446 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U190  ( .ZN(\MAIN/ENGIN/d_d2_stage ), .A(
        \MAIN/ENGIN/STEP_D/n3400 ), .B(\MAIN/ENGIN/STEP_D/n3401 ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_D/U197  ( .ZN(\MAIN/ENGIN/d_exectl_st ), .A(
        \MAIN/ENGIN/STEP_D/n3412 ), .B(\MAIN/ENGIN/STEP_D/n3400 ), .C(
        \MAIN/ENGIN/STEP_D/n3410 ) );
    snl_ao112x1 \MAIN/ENGIN/STEP_D/U203  ( .Z(\MAIN/ENGIN/a_dec_start ), .A(
        \MAIN/ENGIN/STEP_D/n3424 ), .B(\MAIN/ENGIN/STEP_D/n3425 ), .C(
        \MAIN/ENGIN/STEP_D/n3410 ), .D(\MAIN/ENGIN/STEP_D/cst[2] ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_D/U224  ( .ZN(\MAIN/ENGIN/STEP_D/n3437 ), 
        .A(\MAIN/ENGIN/d_cf_stage ), .B(\MAIN/ENGIN/STEP_D/n3412 ), .C(
        pgiaendp) );
    snl_aoi112x0 \MAIN/ENGIN/STEP_D/U199  ( .ZN(
        \MAIN/ENGIN/STEP_D/dec_st2_rst ), .A(\MAIN/ENGIN/STEP_D/n3412 ), .B(
        \MAIN/ENGIN/STEP_D/n3422 ), .C(\MAIN/ENGIN/STEP_D/n3419 ), .D(
        \MAIN/ENGIN/STEP_D/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U202  ( .ZN(ph_dec_dh), .A(
        \MAIN/ENGIN/d_dec_stage ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U210  ( .ZN(\MAIN/ENGIN/STEP_D/n3424 ), .A(
        \MAIN/ENGIN/STEP_D/cst[1] ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U242  ( .ZN(\MAIN/ENGIN/d_step_end ), .A(
        \MAIN/ENGIN/STEP_D/n3414 ) );
    snl_ao022x1 \MAIN/ENGIN/STEP_D/U259  ( .Z(\MAIN/ENGIN/STEP_D/n3445 ), .A(
        \MAIN/exe_end ), .B(\MAIN/ENGIN/STEP_D/cst[2] ), .C(
        \MAIN/ENGIN/STEP_D/n3439 ), .D(\MAIN/ENGIN/STEP_D/n3400 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_D/cst_reg[0]  ( .Q(\MAIN/ENGIN/STEP_D/cst[0] 
        ), .D(\MAIN/ENGIN/STEP_D/tmp2[0] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U237  ( .ZN(\MAIN/ENGIN/STEP_D/n3420 ), .A(
        \MAIN/ENGIN/STEP_D/n3430 ), .B(\MAIN/ENGIN/STEP_D/n3406 ) );
    snl_and34x0 \MAIN/ENGIN/STEP_D/U205  ( .Z(\MAIN/ENGIN/STEP_D/n3426 ), .A(
        \MAIN/ENGIN/STEP_D/cst[1] ), .B(\MAIN/ENGIN/STEP_D/cst[0] ), .C(
        \MAIN/ENGIN/STEP_D/n3427 ), .D(\MAIN/POL_STH ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U219  ( .ZN(\MAIN/ENGIN/STEP_D/n3412 ), .A(
        \MAIN/ENGIN/STEP_D/n3416 ), .B(\MAIN/WP_PC ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U225  ( .ZN(\MAIN/ENGIN/STEP_D/n3438 ), 
        .A(\MAIN/ENGIN/STEP_D/cst[2] ), .B(\MAIN/ENGIN/STEP_D/n3424 ) );
    snl_aoi012x1 \MAIN/ENGIN/STEP_D/U250  ( .ZN(\MAIN/ENGIN/STEP_D/n3446 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/c_decctl_st ), .C(
        \MAIN/ENGIN/STEP_D/n3429 ) );
    snl_ao01b2x0 \MAIN/ENGIN/STEP_D/U222  ( .Z(\MAIN/ENGIN/STEP_D/n3411 ), .A(
        \MAIN/ENGIN/STEP_D/n3434 ), .B(\MAIN/ENGIN/STEP_D/n3435 ), .C(
        \MAIN/ENGIN/status_wr4 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U239  ( .ZN(\MAIN/ENGIN/D_INIT_STAGE ), .A(
        \MAIN/ENGIN/STEP_D/n3435 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U257  ( .ZN(\MAIN/ENGIN/STEP_D/n3440 ), 
        .A(\MAIN/sw_end ), .B(\MAIN/ENGIN/STEP_D/n3413 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U217  ( .ZN(\MAIN/ENGIN/STEP_D/n3427 ), .A(
        \MAIN/ENGIN/STEP_D/cst[3] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U230  ( .ZN(\MAIN/ENGIN/STEP_D/n3410 ), .A(
        \MAIN/ENGIN/STEP_D/n3422 ), .B(\MAIN/ENGIN/STEP_D/n3419 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U245  ( .ZN(\MAIN/ENGIN/STEP_D/n3444 ), .A(
        \MAIN/ENGIN/STEP_D/n3412 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_D/cst_reg[2]  ( .Q(\MAIN/ENGIN/STEP_D/cst[2] 
        ), .D(\MAIN/ENGIN/STEP_D/tmp2[2] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_D/exec_stage_reg  ( .Q(\MAIN/d_exec_stage ), 
        .D(\MAIN/ENGIN/STEP_D/exec_stage278 ), .RN(\MAIN/ENGIN/n3591 ), .CP(
        SCLK) );
    snl_and34x0 \MAIN/ENGIN/STEP_D/U192  ( .Z(\MAIN/ENGIN/STEP_D/n3404 ), .A(
        \MAIN/ENGIN/STEP_D/n3406 ), .B(\MAIN/ENGIN/STEP_D/n3407 ), .C(step4_cf
        ), .D(\MAIN/ENGIN/STEP_D/n3405 ) );
    snl_aoi013x0 \MAIN/ENGIN/STEP_D/U207  ( .ZN(\MAIN/ENGIN/STEP_D/n3417 ), 
        .A(\MAIN/ENGIN/STEP_D/n3412 ), .B(\MAIN/ENGIN/STEP_D/n3429 ), .C(
        \MAIN/ENGIN/STEP_D/n3430 ), .D(step4_cf) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U220  ( .ZN(\MAIN/ENGIN/STEP_D/n3413 ), .A(
        \MAIN/ENGIN/c_decctl_st ) );
    snl_oai233x0 \MAIN/ENGIN/STEP_D/U255  ( .ZN(\MAIN/ENGIN/STEP_D/n3442 ), 
        .A(\MAIN/ENGIN/STEP_D/n3427 ), .B(\MAIN/ENGIN/D_PED4_BR ), .C(
        \MAIN/ENGIN/STEP_D/n3429 ), .D(\MAIN/ENGIN/STEP_D/n3418 ), .E(
        \MAIN/ENGIN/STEP_D/cst[2] ), .F(\MAIN/ENGIN/STEP_D/n3424 ), .G(
        \MAIN/ENGIN/STEP_D/n3428 ), .H(\MAIN/ENGIN/STEP_D/n3436 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_D/cst_reg[3]  ( .Q(\MAIN/ENGIN/STEP_D/cst[3] 
        ), .D(\MAIN/ENGIN/STEP_D/nst[3] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_D/U193  ( .ZN(\MAIN/ENGIN/STEP_D/n3408 ), 
        .A(\MAIN/ENGIN/STEP_D/cst[2] ), .B(\MAIN/ENGIN/STEP_D/n3409 ), .C(
        \MAIN/ENGIN/STEP_D/n3410 ), .D(\MAIN/ENGIN/STEP_D/n3411 ) );
    snl_ao023x1 \MAIN/ENGIN/STEP_D/U194  ( .Z(\MAIN/ENGIN/STEP_D/nst[3] ), .A(
        \MAIN/ENGIN/STEP_D/n3412 ), .B(\MAIN/ENGIN/STEP_D/n3401 ), .C(
        \MAIN/ENGIN/STEP_D/cst[3] ), .D(\MAIN/ENGIN/STEP_D/cf_st2_rst ), .E(
        pgperrh) );
    snl_oai022x1 \MAIN/ENGIN/STEP_D/U195  ( .ZN(\MAIN/ENGIN/d_cfctl_st ), .A(
        \MAIN/ENGIN/STEP_D/n3413 ), .B(\MAIN/ENGIN/STEP_D/n3414 ), .C(
        \MAIN/ENGIN/STEP_D/n3415 ), .D(\MAIN/ENGIN/STEP_D/n3416 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U212  ( .ZN(\MAIN/ENGIN/STEP_D/n3422 ), .A(
        \MAIN/dec_end ) );
    snl_nand03x0 \MAIN/ENGIN/STEP_D/U215  ( .ZN(\MAIN/ENGIN/STEP_D/n3434 ), 
        .A(\MAIN/ENGIN/STEP_D/n3413 ), .B(\MAIN/ENGIN/STEP_D/n3416 ), .C(
        \MAIN/POL_STH ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U229  ( .ZN(\MAIN/ENGIN/STEP_D/n3418 ), .A(
        \MAIN/ENGIN/d_dec_start ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_D/decode_stage_reg  ( .Q(
        \MAIN/ENGIN/d_dec_stage ), .D(\MAIN/ENGIN/STEP_D/decode_stage272 ), 
        .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK) );
    snl_nor03x0 \MAIN/ENGIN/STEP_D/U247  ( .ZN(\MAIN/ENGIN/STEP_D/n3406 ), .A(
        \MAIN/ENGIN/STEP_D/n3424 ), .B(pol_status), .C(
        \MAIN/ENGIN/STEP_D/n3400 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U232  ( .ZN(\MAIN/ENGIN/STEP_D/n3401 ), 
        .A(\MAIN/ENGIN/STEP_D/cst[1] ), .B(\MAIN/ENGIN/STEP_D/n3429 ) );
    snl_aoi123x0 \MAIN/ENGIN/STEP_D/U235  ( .ZN(\MAIN/ENGIN/STEP_D/n3403 ), 
        .A(\MAIN/ENGIN/STEP_D/cst[2] ), .B(\MAIN/ENGIN/STEP_D/cst[1] ), .C(
        pol_status), .D(\MAIN/ENGIN/STEP_D/sw_stage ), .E(
        \MAIN/ENGIN/STEP_D/n3440 ), .F(\MAIN/ENGIN/STEP_D/n3407 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U240  ( .ZN(\MAIN/ENGIN/d_cf_stage ), .A(
        \MAIN/ENGIN/STEP_D/n3436 ) );
    snl_nor03x0 \MAIN/ENGIN/STEP_D/U200  ( .ZN(
        \MAIN/ENGIN/STEP_D/exec_stage278 ), .A(\MAIN/ENGIN/STEP_D/n3423 ), .B(
        \MAIN/ENGIN/STEP_D/n3408 ), .C(\MAIN/ENGIN/STEP_D/n3404 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U209  ( .ZN(\MAIN/ENGIN/STEP_D/n3429 ), .A(
        \MAIN/ENGIN/STEP_D/cst[0] ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U227  ( .ZN(\MAIN/ENGIN/STEP_D/d3_stage ), 
        .A(\MAIN/ENGIN/STEP_D/n3438 ), .B(\MAIN/ENGIN/STEP_D/cst[0] ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U249  ( .ZN(\MAIN/ENGIN/STEP_D/n3425 ), .A(
        \MAIN/ENGIN/STEP_D/n3432 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U252  ( .ZN(\MAIN/ENGIN/STEP_D/tmp2[2] ), 
        .A(\MAIN/ENGIN/STEP_D/n3408 ) );
    snl_ffqrnx1 \MAIN/ENGIN/STEP_D/cst_reg[1]  ( .Q(\MAIN/ENGIN/STEP_D/cst[1] 
        ), .D(\MAIN/ENGIN/STEP_D/tmp2[1] ), .RN(\MAIN/ENGIN/n3591 ), .CP(SCLK)
         );
    snl_invx05 \MAIN/ENGIN/STEP_D/U201  ( .ZN(ph_exe_dh), .A(
        \MAIN/d_exec_stage ) );
    snl_aoi0b12x0 \MAIN/ENGIN/STEP_D/U208  ( .ZN(\MAIN/ENGIN/STEP_D/n3415 ), 
        .A(\MAIN/ENGIN/STEP_D/d3_stage ), .B(\MAIN/ENGIN/c_decctl_st ), .C(
        \MAIN/ENGIN/STEP_D/n3431 ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U213  ( .ZN(\MAIN/ENGIN/STEP_D/n3432 ), 
        .A(\MAIN/ENGIN/STEP_D/n3427 ), .B(\MAIN/ENGIN/STEP_D/n3429 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U234  ( .ZN(\MAIN/ENGIN/STEP_D/n3439 ), .A(
        \MAIN/dec_end ), .B(\MAIN/ENGIN/STEP_D/n3412 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U241  ( .ZN(\MAIN/ENGIN/status_wr4 ), .A(
        \MAIN/ENGIN/STEP_D/n3427 ), .B(\MAIN/ENGIN/STEP_D/n3424 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U226  ( .ZN(\MAIN/ENGIN/STEP_D/sw_stage ), 
        .A(\MAIN/ENGIN/STEP_D/n3438 ), .B(\MAIN/ENGIN/STEP_D/n3429 ) );
    snl_and23x0 \MAIN/ENGIN/STEP_D/U206  ( .Z(\MAIN/ENGIN/STEP_D/n3428 ), .A(
        \MAIN/ENGIN/d_dec_start ), .B(pgperrh), .C(pgiaendp) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U248  ( .ZN(\MAIN/ENGIN/STEP_D/n3443 ), .A(
        \MAIN/ENGIN/STEP_D/n3438 ) );
    snl_oai012x1 \MAIN/ENGIN/STEP_D/U253  ( .ZN(\MAIN/ENGIN/STEP_D/n3405 ), 
        .A(\MAIN/ENGIN/STEP_D/n3426 ), .B(\MAIN/ENGIN/STEP_D/n3430 ), .C(
        \MAIN/ENGIN/STEP_D/n3412 ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U254  ( .ZN(\MAIN/ENGIN/STEP_D/tmp2[1] ), 
        .A(\MAIN/ENGIN/STEP_D/n3404 ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U214  ( .ZN(\MAIN/ENGIN/STEP_D/n3433 ), .A(
        \MAIN/ENGIN/STEP_D/cst[1] ), .B(\MAIN/ENGIN/STEP_D/cst[2] ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/U221  ( .ZN(\MAIN/ENGIN/STEP_D/n3400 ), .A(
        \MAIN/ENGIN/STEP_D/cst[2] ) );
    snl_nand02x1 \MAIN/ENGIN/STEP_D/U233  ( .ZN(\MAIN/ENGIN/STEP_D/n3414 ), 
        .A(\MAIN/ENGIN/STEP_D/sw_stage ), .B(\MAIN/sw_end ) );
    snl_nor02x1 \MAIN/ENGIN/STEP_D/U246  ( .ZN(\MAIN/ENGIN/STEP_D/n3407 ), .A(
        \MAIN/ENGIN/STEP_D/n3445 ), .B(\MAIN/ENGIN/STEP_D/n3419 ) );
    snl_aoi023x0 \MAIN/ENGIN/STEP_D/U228  ( .ZN(\MAIN/ENGIN/STEP_D/n3431 ), 
        .A(\MAIN/ENGIN/c_decctl_st ), .B(\MAIN/ENGIN/STEP_D/n3424 ), .C(
        \MAIN/ENGIN/STEP_D/n3425 ), .D(\MAIN/ENGIN/STEP_D/d3_stage ), .E(
        \MAIN/WP_PC ) );
    snl_and04x1 \CONS/phinc20_1/inc4_1/U7  ( .Z(\CONS/phinc20_1/gp_out[0] ), 
        .A(\pk_saco_lh[7] ), .B(\pk_saco_lh[4] ), .C(\pk_saco_lh[5] ), .D(
        \pk_saco_lh[6] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_1/U8  ( .ZN(\CONS/phinc20_1/inc4_1/n325 
        ), .A(\pk_saco_lh[4] ), .B(1'b1) );
    snl_xor2x0 \CONS/phinc20_1/inc4_1/U13  ( .Z(\CONS/SACO[0] ), .A(
        \pk_saco_lh[4] ), .B(1'b1) );
    snl_nand02x1 \CONS/phinc20_1/inc4_1/U14  ( .ZN(
        \CONS/phinc20_1/inc4_1/n327 ), .A(\pk_saco_lh[6] ), .B(
        \CONS/phinc20_1/inc4_1/n326 ) );
    snl_and12x1 \CONS/phinc20_1/inc4_1/U9  ( .Z(\CONS/phinc20_1/inc4_1/n326 ), 
        .A(\CONS/phinc20_1/inc4_1/n325 ), .B(\pk_saco_lh[5] ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_1/U12  ( .ZN(\CONS/SACO[1] ), .A(
        \pk_saco_lh[5] ), .B(\CONS/phinc20_1/inc4_1/n325 ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_1/U10  ( .ZN(\CONS/SACO[3] ), .A(
        \pk_saco_lh[7] ), .B(\CONS/phinc20_1/inc4_1/n327 ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_1/U11  ( .Z(\CONS/SACO[2] ), .A(
        \pk_saco_lh[6] ), .B(\CONS/phinc20_1/inc4_1/n326 ) );
    snl_and04x1 \CONS/phinc20_1/inc4_2/U7  ( .Z(\CONS/phinc20_1/gp_out[1] ), 
        .A(\pk_saco_lh[11] ), .B(\pk_saco_lh[8] ), .C(\pk_saco_lh[9] ), .D(
        \pk_saco_lh[10] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_2/U8  ( .ZN(\CONS/phinc20_1/inc4_2/n322 
        ), .A(\pk_saco_lh[8] ), .B(\CONS/phinc20_1/gp_out[0] ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_2/U13  ( .Z(\CONS/SACO[4] ), .A(
        \pk_saco_lh[8] ), .B(\CONS/phinc20_1/gp_out[0] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_2/U14  ( .ZN(
        \CONS/phinc20_1/inc4_2/n324 ), .A(\pk_saco_lh[10] ), .B(
        \CONS/phinc20_1/inc4_2/n323 ) );
    snl_and12x1 \CONS/phinc20_1/inc4_2/U9  ( .Z(\CONS/phinc20_1/inc4_2/n323 ), 
        .A(\CONS/phinc20_1/inc4_2/n322 ), .B(\pk_saco_lh[9] ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_2/U12  ( .ZN(\CONS/SACO[5] ), .A(
        \pk_saco_lh[9] ), .B(\CONS/phinc20_1/inc4_2/n322 ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_2/U10  ( .ZN(\CONS/SACO[7] ), .A(
        \pk_saco_lh[11] ), .B(\CONS/phinc20_1/inc4_2/n324 ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_2/U11  ( .Z(\CONS/SACO[6] ), .A(
        \pk_saco_lh[10] ), .B(\CONS/phinc20_1/inc4_2/n323 ) );
    snl_and04x1 \CONS/phinc20_1/inc4_3/U7  ( .Z(\CONS/phinc20_1/gp_out[2] ), 
        .A(\pk_saco_lh[15] ), .B(\pk_saco_lh[12] ), .C(\pk_saco_lh[13] ), .D(
        \pk_saco_lh[14] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_3/U8  ( .ZN(\CONS/phinc20_1/inc4_3/n319 
        ), .A(\pk_saco_lh[12] ), .B(\CONS/phinc20_1/gg_out[1] ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_3/U13  ( .Z(\CONS/SACO[8] ), .A(
        \pk_saco_lh[12] ), .B(\CONS/phinc20_1/gg_out[1] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_3/U14  ( .ZN(
        \CONS/phinc20_1/inc4_3/n321 ), .A(\pk_saco_lh[14] ), .B(
        \CONS/phinc20_1/inc4_3/n320 ) );
    snl_and12x1 \CONS/phinc20_1/inc4_3/U9  ( .Z(\CONS/phinc20_1/inc4_3/n320 ), 
        .A(\CONS/phinc20_1/inc4_3/n319 ), .B(\pk_saco_lh[13] ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_3/U12  ( .ZN(\CONS/SACO[9] ), .A(
        \pk_saco_lh[13] ), .B(\CONS/phinc20_1/inc4_3/n319 ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_3/U10  ( .ZN(\CONS/SACO[11] ), .A(
        \pk_saco_lh[15] ), .B(\CONS/phinc20_1/inc4_3/n321 ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_3/U11  ( .Z(\CONS/SACO[10] ), .A(
        \pk_saco_lh[14] ), .B(\CONS/phinc20_1/inc4_3/n320 ) );
    snl_and04x1 \CONS/phinc20_1/inc4_4/U7  ( .Z(\CONS/phinc20_1/gp_out[3] ), 
        .A(\pk_saco_lh[19] ), .B(\pk_saco_lh[16] ), .C(\pk_saco_lh[17] ), .D(
        \pk_saco_lh[18] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_4/U8  ( .ZN(\CONS/phinc20_1/inc4_4/n316 
        ), .A(\pk_saco_lh[16] ), .B(\CONS/phinc20_1/gg_out[2] ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_4/U13  ( .Z(\CONS/SACO[12] ), .A(
        \pk_saco_lh[16] ), .B(\CONS/phinc20_1/gg_out[2] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_4/U14  ( .ZN(
        \CONS/phinc20_1/inc4_4/n318 ), .A(\pk_saco_lh[18] ), .B(
        \CONS/phinc20_1/inc4_4/n317 ) );
    snl_and12x1 \CONS/phinc20_1/inc4_4/U9  ( .Z(\CONS/phinc20_1/inc4_4/n317 ), 
        .A(\CONS/phinc20_1/inc4_4/n316 ), .B(\pk_saco_lh[17] ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_4/U12  ( .ZN(\CONS/SACO[13] ), .A(
        \pk_saco_lh[17] ), .B(\CONS/phinc20_1/inc4_4/n316 ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_4/U10  ( .ZN(\CONS/SACO[15] ), .A(
        \pk_saco_lh[19] ), .B(\CONS/phinc20_1/inc4_4/n318 ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_4/U11  ( .Z(\CONS/SACO[14] ), .A(
        \pk_saco_lh[18] ), .B(\CONS/phinc20_1/inc4_4/n317 ) );
    snl_and04x1 \CONS/phinc20_1/inc4_5/U7  ( .Z(\CONS/phinc20_1/inc4_5/gp_out 
        ), .A(\pk_saco_lh[23] ), .B(\pk_saco_lh[20] ), .C(\pk_saco_lh[21] ), 
        .D(\pk_saco_lh[22] ) );
    snl_nand02x1 \CONS/phinc20_1/inc4_5/U8  ( .ZN(\CONS/phinc20_1/inc4_5/n311 
        ), .A(\pk_saco_lh[20] ), .B(\CONS/phinc20_1/gg_out[3] ) );
    snl_aoi022x1 \CONS/phinc20_1/inc4_5/U13  ( .ZN(\CONS/SACO[17] ), .A(
        \pk_saco_lh[21] ), .B(\CONS/phinc20_1/inc4_5/n315 ), .C(
        \CONS/phinc20_1/inc4_5/n312 ), .D(\CONS/phinc20_1/inc4_5/n311 ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_5/U14  ( .Z(\CONS/SACO[16] ), .A(
        \pk_saco_lh[20] ), .B(\CONS/phinc20_1/gg_out[3] ) );
    snl_invx05 \CONS/phinc20_1/inc4_5/U9  ( .ZN(\CONS/phinc20_1/inc4_5/n312 ), 
        .A(\pk_saco_lh[21] ) );
    snl_xor2x0 \CONS/phinc20_1/inc4_5/U12  ( .Z(\CONS/SACO[18] ), .A(
        \pk_saco_lh[22] ), .B(\CONS/phinc20_1/inc4_5/n313 ) );
    snl_nor02x1 \CONS/phinc20_1/inc4_5/U10  ( .ZN(\CONS/phinc20_1/inc4_5/n313 
        ), .A(\CONS/phinc20_1/inc4_5/n312 ), .B(\CONS/phinc20_1/inc4_5/n311 )
         );
    snl_nand02x1 \CONS/phinc20_1/inc4_5/U15  ( .ZN(
        \CONS/phinc20_1/inc4_5/n314 ), .A(\pk_saco_lh[22] ), .B(
        \CONS/phinc20_1/inc4_5/n313 ) );
    snl_xnor2x0 \CONS/phinc20_1/inc4_5/U11  ( .ZN(\CONS/SACO[19] ), .A(
        \pk_saco_lh[23] ), .B(\CONS/phinc20_1/inc4_5/n314 ) );
    snl_invx05 \CONS/phinc20_1/inc4_5/U16  ( .ZN(\CONS/phinc20_1/inc4_5/n315 ), 
        .A(\CONS/phinc20_1/inc4_5/n311 ) );
    snl_and04x1 \CODEIF/inc19_1/inc4_1/U7  ( .Z(\CODEIF/inc19_1/gp_out[0] ), 
        .A(\CODEIF/pfctr[3] ), .B(\CODEIF/pfctr[0] ), .C(\CODEIF/pfctr[1] ), 
        .D(\CODEIF/pfctr[2] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_1/U8  ( .ZN(
        \CODEIF/inc19_1/inc4_1/n3760 ), .A(\CODEIF/pfctr[0] ), .B(1'b1) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_1/U13  ( .Z(\CODEIF/pgctrinc[0] ), .A(
        \CODEIF/pfctr[0] ), .B(1'b1) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_1/U14  ( .ZN(
        \CODEIF/inc19_1/inc4_1/n3762 ), .A(\CODEIF/pfctr[2] ), .B(
        \CODEIF/inc19_1/inc4_1/n3761 ) );
    snl_and12x1 \CODEIF/inc19_1/inc4_1/U9  ( .Z(\CODEIF/inc19_1/inc4_1/n3761 ), 
        .A(\CODEIF/inc19_1/inc4_1/n3760 ), .B(\CODEIF/pfctr[1] ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_1/U12  ( .ZN(\CODEIF/pgctrinc[1] ), .A(
        \CODEIF/pfctr[1] ), .B(\CODEIF/inc19_1/inc4_1/n3760 ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_1/U10  ( .ZN(\CODEIF/pgctrinc[3] ), .A(
        \CODEIF/pfctr[3] ), .B(\CODEIF/inc19_1/inc4_1/n3762 ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_1/U11  ( .Z(\CODEIF/pgctrinc[2] ), .A(
        \CODEIF/pfctr[2] ), .B(\CODEIF/inc19_1/inc4_1/n3761 ) );
    snl_and04x1 \CODEIF/inc19_1/inc4_2/U7  ( .Z(\CODEIF/inc19_1/gp_out[1] ), 
        .A(\CODEIF/pfctr[7] ), .B(\CODEIF/pfctr[4] ), .C(\CODEIF/pfctr[5] ), 
        .D(\CODEIF/pfctr[6] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_2/U8  ( .ZN(
        \CODEIF/inc19_1/inc4_2/n3757 ), .A(\CODEIF/pfctr[4] ), .B(
        \CODEIF/inc19_1/gp_out[0] ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_2/U13  ( .Z(\CODEIF/pgctrinc[4] ), .A(
        \CODEIF/pfctr[4] ), .B(\CODEIF/inc19_1/gp_out[0] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_2/U14  ( .ZN(
        \CODEIF/inc19_1/inc4_2/n3759 ), .A(\CODEIF/pfctr[6] ), .B(
        \CODEIF/inc19_1/inc4_2/n3758 ) );
    snl_and12x1 \CODEIF/inc19_1/inc4_2/U9  ( .Z(\CODEIF/inc19_1/inc4_2/n3758 ), 
        .A(\CODEIF/inc19_1/inc4_2/n3757 ), .B(\CODEIF/pfctr[5] ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_2/U12  ( .ZN(\CODEIF/pgctrinc[5] ), .A(
        \CODEIF/pfctr[5] ), .B(\CODEIF/inc19_1/inc4_2/n3757 ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_2/U10  ( .ZN(\CODEIF/pgctrinc[7] ), .A(
        \CODEIF/pfctr[7] ), .B(\CODEIF/inc19_1/inc4_2/n3759 ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_2/U11  ( .Z(\CODEIF/pgctrinc[6] ), .A(
        \CODEIF/pfctr[6] ), .B(\CODEIF/inc19_1/inc4_2/n3758 ) );
    snl_and04x1 \CODEIF/inc19_1/inc4_3/U7  ( .Z(\CODEIF/inc19_1/gp_out[2] ), 
        .A(\CODEIF/pfctr[11] ), .B(\CODEIF/pfctr[8] ), .C(\CODEIF/pfctr[9] ), 
        .D(\CODEIF/pfctr[10] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_3/U8  ( .ZN(
        \CODEIF/inc19_1/inc4_3/n3656 ), .A(\CODEIF/pfctr[8] ), .B(
        \CODEIF/inc19_1/gg_out[1] ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_3/U13  ( .Z(\CODEIF/pgctrinc[8] ), .A(
        \CODEIF/pfctr[8] ), .B(\CODEIF/inc19_1/gg_out[1] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_3/U14  ( .ZN(
        \CODEIF/inc19_1/inc4_3/n3756 ), .A(\CODEIF/pfctr[10] ), .B(
        \CODEIF/inc19_1/inc4_3/n3755 ) );
    snl_and12x1 \CODEIF/inc19_1/inc4_3/U9  ( .Z(\CODEIF/inc19_1/inc4_3/n3755 ), 
        .A(\CODEIF/inc19_1/inc4_3/n3656 ), .B(\CODEIF/pfctr[9] ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_3/U12  ( .ZN(\CODEIF/pgctrinc[9] ), .A(
        \CODEIF/pfctr[9] ), .B(\CODEIF/inc19_1/inc4_3/n3656 ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_3/U10  ( .ZN(\CODEIF/pgctrinc[11] ), .A(
        \CODEIF/pfctr[11] ), .B(\CODEIF/inc19_1/inc4_3/n3756 ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_3/U11  ( .Z(\CODEIF/pgctrinc[10] ), .A(
        \CODEIF/pfctr[10] ), .B(\CODEIF/inc19_1/inc4_3/n3755 ) );
    snl_and04x1 \CODEIF/inc19_1/inc4_4/U7  ( .Z(\CODEIF/inc19_1/gp_out[3] ), 
        .A(\CODEIF/pfctr[15] ), .B(\CODEIF/pfctr[12] ), .C(\CODEIF/pfctr[13] ), 
        .D(\CODEIF/pfctr[14] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_4/U8  ( .ZN(
        \CODEIF/inc19_1/inc4_4/n3650 ), .A(\CODEIF/pfctr[12] ), .B(
        \CODEIF/inc19_1/gg_out[2] ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_4/U13  ( .Z(\CODEIF/pgctrinc[12] ), .A(
        \CODEIF/pfctr[12] ), .B(\CODEIF/inc19_1/gg_out[2] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_4/U14  ( .ZN(
        \CODEIF/inc19_1/inc4_4/n3654 ), .A(\CODEIF/pfctr[14] ), .B(
        \CODEIF/inc19_1/inc4_4/n3652 ) );
    snl_and12x1 \CODEIF/inc19_1/inc4_4/U9  ( .Z(\CODEIF/inc19_1/inc4_4/n3652 ), 
        .A(\CODEIF/inc19_1/inc4_4/n3650 ), .B(\CODEIF/pfctr[13] ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_4/U12  ( .ZN(\CODEIF/pgctrinc[13] ), .A(
        \CODEIF/pfctr[13] ), .B(\CODEIF/inc19_1/inc4_4/n3650 ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_4/U10  ( .ZN(\CODEIF/inc19_1/n3763 ), .A(
        \CODEIF/pfctr[15] ), .B(\CODEIF/inc19_1/inc4_4/n3654 ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_4/U11  ( .Z(\CODEIF/pgctrinc[14] ), .A(
        \CODEIF/pfctr[14] ), .B(\CODEIF/inc19_1/inc4_4/n3652 ) );
    snl_and04x1 \CODEIF/inc19_1/inc4_5/U7  ( .Z(\CODEIF/inc19_1/inc4_5/gp_out 
        ), .A(\CODEIF/pfctr[18] ), .B(\CODEIF/pfctr[15] ), .C(
        \CODEIF/pfctr[16] ), .D(\CODEIF/pfctr[17] ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_5/U8  ( .ZN(
        \CODEIF/inc19_1/inc4_5/n3640 ), .A(\CODEIF/pfctr[15] ), .B(
        \CODEIF/inc19_1/gg_out[3] ) );
    snl_aoi022x1 \CODEIF/inc19_1/inc4_5/U13  ( .ZN(\CODEIF/pgctrinc[16] ), .A(
        \CODEIF/pfctr[16] ), .B(\CODEIF/inc19_1/inc4_5/n3648 ), .C(
        \CODEIF/inc19_1/inc4_5/n3642 ), .D(\CODEIF/inc19_1/inc4_5/n3640 ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_5/U14  ( .Z(\CODEIF/inc19_1/n3764 ), .A(
        \CODEIF/pfctr[15] ), .B(\CODEIF/inc19_1/gg_out[3] ) );
    snl_invx05 \CODEIF/inc19_1/inc4_5/U9  ( .ZN(\CODEIF/inc19_1/inc4_5/n3642 ), 
        .A(\CODEIF/pfctr[16] ) );
    snl_xor2x0 \CODEIF/inc19_1/inc4_5/U12  ( .Z(\CODEIF/pgctrinc[17] ), .A(
        \CODEIF/pfctr[17] ), .B(\CODEIF/inc19_1/inc4_5/n3644 ) );
    snl_nor02x1 \CODEIF/inc19_1/inc4_5/U10  ( .ZN(
        \CODEIF/inc19_1/inc4_5/n3644 ), .A(\CODEIF/inc19_1/inc4_5/n3642 ), .B(
        \CODEIF/inc19_1/inc4_5/n3640 ) );
    snl_nand02x1 \CODEIF/inc19_1/inc4_5/U15  ( .ZN(
        \CODEIF/inc19_1/inc4_5/n3646 ), .A(\CODEIF/pfctr[17] ), .B(
        \CODEIF/inc19_1/inc4_5/n3644 ) );
    snl_xnor2x0 \CODEIF/inc19_1/inc4_5/U11  ( .ZN(\CODEIF/pgctrinc[18] ), .A(
        \CODEIF/pfctr[18] ), .B(\CODEIF/inc19_1/inc4_5/n3646 ) );
    snl_invx05 \CODEIF/inc19_1/inc4_5/U16  ( .ZN(\CODEIF/inc19_1/inc4_5/n3648 
        ), .A(\CODEIF/inc19_1/inc4_5/n3640 ) );
    snl_and08x1 \UPIF/RCTL/regfile_1/U6  ( .Z(\UPIF/RCTL/reg_file_h ), .A(PA
        [29]), .B(PA[27]), .C(\UPIF/RCTL/regfile_1/n1016 ), .D(PA[13]), .E(
        \UPIF/RCTL/regfile_1/n1017 ), .F(\UPIF/RCTL/regfile_1/n1018 ), .G(
        \UPIF/RCTL/regfile_1/n1019 ), .H(\UPIF/RCTL/regfile_1/n1020 ) );
    snl_nor03x0 \UPIF/RCTL/regfile_1/U7  ( .ZN(\UPIF/RCTL/regfile_1/n1019 ), 
        .A(PA[28]), .B(PA[31]), .C(PA[30]) );
    snl_nor03x0 \UPIF/RCTL/regfile_1/U8  ( .ZN(\UPIF/RCTL/regfile_1/n1018 ), 
        .A(PA[24]), .B(PA[26]), .C(PA[25]) );
    snl_nor02x1 \UPIF/RCTL/regfile_1/U13  ( .ZN(\UPIF/RCTL/regfile_1/n1016 ), 
        .A(PA[12]), .B(PA[11]) );
    snl_nor02x1 \UPIF/RCTL/regfile_1/U9  ( .ZN(\UPIF/RCTL/regfile_1/n1021 ), 
        .A(PA[23]), .B(PA[22]) );
    snl_and34x0 \UPIF/RCTL/regfile_1/U12  ( .Z(\UPIF/RCTL/regfile_1/n1017 ), 
        .A(PA[15]), .B(PA[14]), .C(PA[16]), .D(\UPIF/RCTL/regfile_1/n1022 ) );
    snl_and34x0 \UPIF/RCTL/regfile_1/U10  ( .Z(\UPIF/RCTL/regfile_1/n1020 ), 
        .A(PA[20]), .B(PA[19]), .C(PA[21]), .D(\UPIF/RCTL/regfile_1/n1021 ) );
    snl_nor02x1 \UPIF/RCTL/regfile_1/U11  ( .ZN(\UPIF/RCTL/regfile_1/n1022 ), 
        .A(PA[18]), .B(PA[17]) );
    snl_oai013x0 \REGF/pbmemff31/SACNST/U23  ( .ZN(
        \REGF/pbmemff31/SACNST/*cell*5426/U1/CONTROL2 ), .A(
        \REGF/pbmemff31/SACNST/n5645 ), .B(\pk_rwrit_h[48] ), .C(ph_stregwt_h), 
        .D(\REGF/pbmemff31/SACNST/n5646 ) );
    snl_invx05 \REGF/pbmemff31/SACNST/U24  ( .ZN(\REGF/pbmemff31/SACNST/n5645 
        ), .A(\REGF/pbmemff31/DO_SACONS ) );
    snl_oai012x1 \REGF/pbmemff31/SACNST/U25  ( .ZN(
        \REGF/pbmemff31/SACNST/n5646 ), .A(\REGF/pbmemff31/DO_SACONS ), .B(
        ph_sacons_h), .C(ad_latch) );
    snl_ffqrnx1 \REGF/pbmemff31/SACNST/DO_SACONS_reg  ( .Q(
        \REGF/pbmemff31/DO_SACONS ), .D(
        \REGF/pbmemff31/SACNST/*cell*5426/U1/CONTROL2 ), .RN(
        \REGF/pbmemff31/n5648 ), .CP(SCLK) );
    snl_or02x1 \ALUSHT/ALU/dec32/U6  ( .Z(\ALUSHT/ALU/dec32/gcarry[1] ), .A(
        \ALUSHT/ALU/dec32/gg_out[0] ), .B(\ALUSHT/ALU/dec32/gg_out[1] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/U8  ( .ZN(\ALUSHT/ALU/dec32/n1801 ), .A(
        \ALUSHT/ALU/dec32/gg_out[5] ), .B(\ALUSHT/ALU/dec32/gcarry[4] ) );
    snl_invx05 \ALUSHT/ALU/dec32/U12  ( .ZN(\ALUSHT/ALU/dec32/gcarry[5] ), .A(
        \ALUSHT/ALU/dec32/n1801 ) );
    snl_nand12x1 \ALUSHT/ALU/dec32/U9  ( .ZN(\ALUSHT/ALU/dec32/gcarry[6] ), 
        .A(\ALUSHT/ALU/dec32/gg_out[6] ), .B(\ALUSHT/ALU/dec32/n1801 ) );
    snl_or02x1 \ALUSHT/ALU/dec32/U7  ( .Z(\ALUSHT/ALU/dec32/gcarry[4] ), .A(
        \ALUSHT/ALU/dec32/gg_out[4] ), .B(\ALUSHT/ALU/dec32/gcarry[3] ) );
    snl_or02x1 \ALUSHT/ALU/dec32/U10  ( .Z(\ALUSHT/ALU/dec32/gcarry[2] ), .A(
        \ALUSHT/ALU/dec32/gg_out[2] ), .B(\ALUSHT/ALU/dec32/gcarry[1] ) );
    snl_or02x1 \ALUSHT/ALU/dec32/U11  ( .Z(\ALUSHT/ALU/dec32/gcarry[3] ), .A(
        \ALUSHT/ALU/dec32/gg_out[3] ), .B(\ALUSHT/ALU/dec32/gcarry[2] ) );
    snl_xnor2x0 \ALUSHT/ALU/add32/U13  ( .ZN(\ALUSHT/ALU/pkovf32 ), .A(
        \ALUSHT/ALU/add32/c_last ), .B(\ALUSHT/ALU/add32/n1635 ) );
    snl_invx05 \ALUSHT/ALU/add32/U14  ( .ZN(\ALUSHT/ALU/add32/n1390 ), .A(
        \ALUSHT/ALU/add32/gp_out[1] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/U8  ( .ZN(\ALUSHT/ALU/add32/cin_stg[1] ), 
        .A(\ALUSHT/ALU/add32/n1389 ), .B(\ALUSHT/ALU/add32/n1390 ), .C(
        \ALUSHT/ALU/add32/n1394 ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/U12  ( .ZN(\ALUSHT/ALU/add32/n1635 ), .A(
        \ALUSHT/ALU/add32/gp_out[5] ), .B(\ALUSHT/ALU/add32/cin_stg[4] ), .C(
        \ALUSHT/ALU/add32/gg_out[5] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/U9  ( .ZN(\ALUSHT/ALU/add32/n1389 ), .A(
        \ALUSHT/ALU/add32/gp_out[0] ), .B(\ALUSHT/ALU/pkaddcin ), .C(
        \ALUSHT/ALU/add32/gg_out[0] ) );
    snl_ao012x1 \ALUSHT/ALU/add32/U7  ( .Z(\ALUSHT/ALU/add32/cin_stg[3] ), .A(
        \ALUSHT/ALU/add32/gp_out[3] ), .B(\ALUSHT/ALU/add32/cin_stg[2] ), .C(
        \ALUSHT/ALU/add32/gg_out[3] ) );
    snl_ao012x1 \ALUSHT/ALU/add32/U10  ( .Z(\ALUSHT/ALU/add32/cin_stg[4] ), 
        .A(\ALUSHT/ALU/add32/gp_out[4] ), .B(\ALUSHT/ALU/add32/cin_stg[3] ), 
        .C(\ALUSHT/ALU/add32/gg_out[4] ) );
    snl_invx05 \ALUSHT/ALU/add32/U15  ( .ZN(\ALUSHT/ALU/add32/n1394 ), .A(
        \ALUSHT/ALU/add32/gg_out[1] ) );
    snl_ao012x1 \ALUSHT/ALU/add32/U11  ( .Z(\ALUSHT/ALU/add32/cin_stg[2] ), 
        .A(\ALUSHT/ALU/add32/gp_out[2] ), .B(\ALUSHT/ALU/add32/cin_stg[1] ), 
        .C(\ALUSHT/ALU/add32/gg_out[2] ) );
    snl_invx05 \ALUSHT/ALU/add32/U16  ( .ZN(\ALUSHT/ALU/add32/cin_stg[0] ), 
        .A(\ALUSHT/ALU/add32/n1389 ) );
    snl_nor02x1 \ALUSHT/ALU/cmp32/U13  ( .ZN(\ALUSHT/ALU/cmp32/n1218 ), .A(
        \ALUSHT/ALU/cmp32/n1216 ), .B(\ALUSHT/ALU/cmp32/n1219 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/U14  ( .ZN(\ALUSHT/ALU/cmp32/n1214 ), .A(
        \ALUSHT/ALU/cmp32/geqflg[2] ) );
    snl_nand12x1 \ALUSHT/ALU/cmp32/U8  ( .ZN(\ALUSHT/ALU/pkgtflg ), .A(
        \ALUSHT/ALU/cmp32/ggflg[7] ), .B(\ALUSHT/ALU/cmp32/n1211 ) );
    snl_and08x1 \ALUSHT/ALU/cmp32/U7  ( .Z(\ALUSHT/ALU/pkeqflg ), .A(
        \ALUSHT/ALU/cmp32/geqflg[0] ), .B(\ALUSHT/ALU/cmp32/geqflg[7] ), .C(
        \ALUSHT/ALU/cmp32/geqflg[6] ), .D(\ALUSHT/ALU/cmp32/geqflg[5] ), .E(
        \ALUSHT/ALU/cmp32/geqflg[4] ), .F(\ALUSHT/ALU/cmp32/geqflg[3] ), .G(
        \ALUSHT/ALU/cmp32/geqflg[2] ), .H(\ALUSHT/ALU/cmp32/geqflg[1] ) );
    snl_aoi012x1 \ALUSHT/ALU/cmp32/U9  ( .ZN(\ALUSHT/ALU/cmp32/n1212 ), .A(
        \ALUSHT/ALU/cmp32/ggflg[0] ), .B(\ALUSHT/ALU/cmp32/geqflg[1] ), .C(
        \ALUSHT/ALU/cmp32/ggflg[1] ) );
    snl_aoi012x1 \ALUSHT/ALU/cmp32/U12  ( .ZN(\ALUSHT/ALU/cmp32/n1216 ), .A(
        \ALUSHT/ALU/cmp32/geqflg[5] ), .B(\ALUSHT/ALU/cmp32/n1217 ), .C(
        \ALUSHT/ALU/cmp32/ggflg[5] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/U15  ( .ZN(\ALUSHT/ALU/cmp32/n1219 ), .A(
        \ALUSHT/ALU/cmp32/geqflg[6] ) );
    snl_nor02x1 \ALUSHT/ALU/cmp32/U10  ( .ZN(\ALUSHT/ALU/cmp32/n1213 ), .A(
        \ALUSHT/ALU/cmp32/n1212 ), .B(\ALUSHT/ALU/cmp32/n1214 ) );
    snl_nand12x1 \ALUSHT/ALU/cmp32/U17  ( .ZN(\ALUSHT/ALU/cmp32/n1217 ), .A(
        \ALUSHT/ALU/cmp32/ggflg[4] ), .B(\ALUSHT/ALU/cmp32/n1220 ) );
    snl_oa012x1 \ALUSHT/ALU/cmp32/U11  ( .Z(\ALUSHT/ALU/cmp32/n1215 ), .A(
        \ALUSHT/ALU/cmp32/n1213 ), .B(\ALUSHT/ALU/cmp32/ggflg[2] ), .C(
        \ALUSHT/ALU/cmp32/geqflg[3] ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/U16  ( .ZN(\ALUSHT/ALU/cmp32/n1220 ), .A(
        \ALUSHT/ALU/cmp32/n1215 ), .B(\ALUSHT/ALU/cmp32/ggflg[3] ), .C(
        \ALUSHT/ALU/cmp32/geqflg[4] ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/U18  ( .ZN(\ALUSHT/ALU/cmp32/n1211 ), .A(
        \ALUSHT/ALU/cmp32/n1218 ), .B(\ALUSHT/ALU/cmp32/ggflg[6] ), .C(
        \ALUSHT/ALU/cmp32/geqflg[7] ) );
    snl_and02x1 \ALUSHT/ALU/inc32/U6  ( .Z(\ALUSHT/ALU/inc32/gg_out[6] ), .A(
        \ALUSHT/ALU/inc32/gg_out[5] ), .B(\ALUSHT/ALU/inc32/gp_out[6] ) );
    snl_and02x1 \ALUSHT/ALU/inc32/U8  ( .Z(\ALUSHT/ALU/inc32/gg_out[2] ), .A(
        \ALUSHT/ALU/inc32/gp_out[2] ), .B(\ALUSHT/ALU/inc32/gg_out[1] ) );
    snl_and02x1 \ALUSHT/ALU/inc32/U9  ( .Z(\ALUSHT/ALU/inc32/gg_out[3] ), .A(
        \ALUSHT/ALU/inc32/gp_out[3] ), .B(\ALUSHT/ALU/inc32/gg_out[2] ) );
    snl_and02x1 \ALUSHT/ALU/inc32/U7  ( .Z(\ALUSHT/ALU/inc32/gg_out[1] ), .A(
        \ALUSHT/ALU/inc32/gp_out[1] ), .B(\ALUSHT/ALU/inc32/gp_out[0] ) );
    snl_and02x1 \ALUSHT/ALU/inc32/U10  ( .Z(\ALUSHT/ALU/inc32/gg_out[4] ), .A(
        \ALUSHT/ALU/inc32/gp_out[4] ), .B(\ALUSHT/ALU/inc32/gg_out[3] ) );
    snl_and02x1 \ALUSHT/ALU/inc32/U11  ( .Z(\ALUSHT/ALU/inc32/gg_out[5] ), .A(
        \ALUSHT/ALU/inc32/gp_out[5] ), .B(\ALUSHT/ALU/inc32/gg_out[4] ) );
    snl_oai112x0 \MAIN/STM/SEQMG/U112  ( .ZN(lbus_locken_h), .A(
        \MAIN/STM/seq_end ), .B(\MAIN/STM/SEQMG/n3345 ), .C(
        \MAIN/STM/SEQMG/n3346 ), .D(\MAIN/STM/SEQMG/n3347 ) );
    snl_nand12x1 \MAIN/STM/SEQMG/U113  ( .ZN(\MAIN/STM/srgfilewren_h ), .A(
        \MAIN/STM/exec_eoc ), .B(\MAIN/STM/SEQMG/n3348 ) );
    snl_nor03x0 \MAIN/STM/SEQMG/U114  ( .ZN(\MAIN/STM/exe_1st ), .A(
        \MAIN/STM/SEQMG/n3349 ), .B(\MAIN/single_write ), .C(
        \MAIN/STM/SEQMG/n3347 ) );
    snl_nand02x1 \MAIN/STM/SEQMG/U121  ( .ZN(\MAIN/STM/seq_doing ), .A(
        \MAIN/STM/SEQMG/n3353 ), .B(\MAIN/STM/SEQMG/n3345 ) );
    snl_nor02x1 \MAIN/STM/SEQMG/U126  ( .ZN(\MAIN/STM/SEQMG/n3361 ), .A(
        \MAIN/STM/SEQMG/n3345 ), .B(\MAIN/STM/execute_err ) );
    snl_nand12x1 \MAIN/STM/SEQMG/U134  ( .ZN(\MAIN/STM/SEQMG/n3349 ), .A(
        \MAIN/single_read ), .B(\MAIN/STM/SEQMG/n3351 ) );
    snl_ao022x1 \MAIN/STM/SEQMG/U141  ( .Z(\MAIN/STM/SEQMG/temp[1] ), .A(
        \MAIN/STM/SEQMG/n3362 ), .B(\MAIN/STM/seq_end ), .C(
        \MAIN/STM/SEQMG/eqst[1] ), .D(\MAIN/STM/SEQMG/n3357 ) );
    snl_ffqrnx1 \MAIN/STM/SEQMG/eqst_reg[1]  ( .Q(\MAIN/STM/SEQMG/eqst[1] ), 
        .D(\MAIN/STM/SEQMG/temp[1] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_or02x1 \MAIN/STM/SEQMG/U128  ( .Z(\MAIN/STM/SEQMG/n3360 ), .A(
        \MAIN/ph_rmw1h ), .B(ph_rmw2h) );
    snl_nor02x1 \MAIN/STM/SEQMG/U133  ( .ZN(\MAIN/STM/SEQMG/n3351 ), .A(
        \MAIN/STM/SEQMG/n3360 ), .B(\MAIN/ph_rrmwh ) );
    snl_ao1b1b3x0 \MAIN/STM/SEQMG/U115  ( .Z(\MAIN/STM/SEQMG/n3350 ), .A(
        \MAIN/STM/execute_err ), .B(\MAIN/ADROVH ), .C(\MAIN/STM/SEQMG/n3351 ), 
        .D(\MAIN/STM/SEQMG/n3353 ), .E(\MAIN/STM/SEQMG/n3352 ) );
    snl_oa012x1 \MAIN/STM/SEQMG/U120  ( .Z(ph_lockh), .A(
        \MAIN/STM/SEQMG/temp[1] ), .B(ph_rmw2h), .C(lbus_locken_h) );
    snl_invx05 \MAIN/STM/SEQMG/U132  ( .ZN(\MAIN/STM/SEQMG/n3356 ), .A(
        \MAIN/single_write ) );
    snl_nand03x0 \MAIN/STM/SEQMG/U129  ( .ZN(\MAIN/STM/SEQMG/n3348 ), .A(
        \MAIN/STM/seq_end ), .B(\MAIN/STM/SEQMG/n3353 ), .C(
        \MAIN/STM/SEQMG/n3361 ) );
    snl_invx05 \MAIN/STM/SEQMG/U140  ( .ZN(\MAIN/STM/SEQMG/n3355 ), .A(
        \MAIN/STM/SEQMG/n3349 ) );
    snl_oai023x0 \MAIN/STM/SEQMG/U116  ( .ZN(\MAIN/STM/exe_1st_r ), .A(
        \MAIN/STM/SEQMG/n3348 ), .B(\MAIN/ADROVH ), .C(\MAIN/STM/SEQMG/n3354 ), 
        .D(\MAIN/STM/SEQMG/n3355 ), .E(\MAIN/STM/SEQMG/n3347 ) );
    snl_nor02x1 \MAIN/STM/SEQMG/U117  ( .ZN(\MAIN/STM/exe_1st_w ), .A(
        \MAIN/STM/SEQMG/n3347 ), .B(\MAIN/STM/SEQMG/n3356 ) );
    snl_nor03x0 \MAIN/STM/SEQMG/U119  ( .ZN(\MAIN/ovferlth ), .A(
        \MAIN/STM/SEQMG/n3359 ), .B(\MAIN/STM/SEQMG/n3351 ), .C(
        \MAIN/STM/SEQMG/n3348 ) );
    snl_invx05 \MAIN/STM/SEQMG/U127  ( .ZN(\MAIN/STM/SEQMG/n3354 ), .A(
        \MAIN/ph_rrmwh ) );
    snl_aoi012x1 \MAIN/STM/SEQMG/U135  ( .ZN(\MAIN/STM/SEQMG/n3362 ), .A(
        \MAIN/STM/SEQMG/eqst[1] ), .B(\MAIN/STM/execute_err ), .C(
        \MAIN/STM/SEQMG/n3345 ) );
    snl_nor03x0 \MAIN/STM/SEQMG/U137  ( .ZN(\MAIN/STM/exec_eoc ), .A(
        \MAIN/STM/SEQMG/n3353 ), .B(\MAIN/STM/SEQMG/n3361 ), .C(
        \MAIN/STM/SEQMG/n3357 ) );
    snl_invx05 \MAIN/STM/SEQMG/U142  ( .ZN(\MAIN/STM/exe_2nd ), .A(
        \MAIN/STM/SEQMG/n3350 ) );
    snl_aoi013x0 \MAIN/STM/SEQMG/U122  ( .ZN(\MAIN/STM/SEQMG/n3358 ), .A(
        \MAIN/STM/SEQMG/n3360 ), .B(\MAIN/STM/SEQMG/n3359 ), .C(
        \MAIN/STM/SEQMG/eqst[0] ), .D(ph_ovfihbh) );
    snl_invx05 \MAIN/STM/SEQMG/U125  ( .ZN(\MAIN/STM/SEQMG/n3345 ), .A(
        \MAIN/STM/SEQMG/eqst[0] ) );
    snl_nand04x0 \MAIN/STM/SEQMG/U139  ( .ZN(\MAIN/STM/SEQMG/n3346 ), .A(
        \MAIN/ph_rrmwh ), .B(\MAIN/STM/SEQMG/n3361 ), .C(
        \MAIN/STM/SEQMG/n3353 ), .D(\MAIN/STM/SEQMG/n3359 ) );
    snl_invx05 \MAIN/STM/SEQMG/U123  ( .ZN(\MAIN/STM/SEQMG/n3353 ), .A(
        \MAIN/STM/SEQMG/eqst[1] ) );
    snl_invx05 \MAIN/STM/SEQMG/U130  ( .ZN(\MAIN/STM/SEQMG/n3359 ), .A(
        \MAIN/ADROVH ) );
    snl_nor02x1 \MAIN/STM/SEQMG/U138  ( .ZN(ph_ovfihbh), .A(
        \MAIN/STM/SEQMG/n3345 ), .B(\MAIN/STM/SEQMG/n3353 ) );
    snl_nor03x0 \MAIN/STM/SEQMG/U118  ( .ZN(\MAIN/STM/exe_2nd_w ), .A(
        \MAIN/STM/SEQMG/n3357 ), .B(\MAIN/STM/execute_err ), .C(
        \MAIN/STM/SEQMG/n3358 ) );
    snl_invx05 \MAIN/STM/SEQMG/U124  ( .ZN(\MAIN/STM/SEQMG/n3357 ), .A(
        \MAIN/STM/seq_end ) );
    snl_nand13x1 \MAIN/STM/SEQMG/U131  ( .ZN(\MAIN/STM/SEQMG/n3347 ), .A(
        \MAIN/STM/seq_doing ), .B(\MAIN/seq_enable ), .C(st_exectl) );
    snl_nand02x1 \MAIN/STM/SEQMG/U136  ( .ZN(\MAIN/STM/SEQMG/n3352 ), .A(
        \MAIN/STM/SEQMG/eqst[0] ), .B(\MAIN/STM/seq_end ) );
    snl_sffqrnx1 \MAIN/STM/SEQMG/b_stage_reg  ( .Q(stage_b), .D(lbus_locken_h), 
        .RN(\MAIN/n3611 ), .SD(1'b0), .SE(\MAIN/STM/SEQMG/temp[1] ), .CP(SCLK)
         );
    snl_ffqrnx1 \MAIN/STM/SEQMG/eqst_reg[0]  ( .Q(\MAIN/STM/SEQMG/eqst[0] ), 
        .D(lbus_locken_h), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_ffqrnx1 \MAIN/STM/SEQMG/stage_2_reg  ( .Q(stage_2), .D(
        \MAIN/STM/SEQMG/temp[1] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nor02x1 \MAIN/STM/NS/U31  ( .ZN(\MAIN/STM/exec_eoc1 ), .A(
        \MAIN/STM/seq_doing ), .B(\MAIN/STM/NS/n3338 ) );
    snl_and02x1 \MAIN/STM/NS/U32  ( .Z(\MAIN/STM/exec_end1 ), .A(
        \MAIN/STM/NS/est[1] ), .B(\MAIN/STM/seq_doing ) );
    snl_aoi012x1 \MAIN/STM/NS/U33  ( .ZN(\MAIN/STM/NS/n3339 ), .A(
        \MAIN/STM/NS/n3340 ), .B(\MAIN/STM/NS/n3341 ), .C(\MAIN/STM/NS/est[1] 
        ) );
    snl_oai223x0 \MAIN/STM/NS/U34  ( .ZN(\MAIN/STM/NS/nst[0] ), .A(
        \MAIN/STM/NS/n3342 ), .B(\MAIN/seq_enable ), .C(\MAIN/STM/NS/n3343 ), 
        .D(\MAIN/STM/NS/n3343 ), .E(\MAIN/STM/NS/n3340 ), .F(
        \MAIN/STM/NS/n3339 ), .G(\MAIN/STM/NS/n3344 ) );
    snl_invx05 \MAIN/STM/NS/U35  ( .ZN(\MAIN/STM/NS/n3344 ), .A(
        \MAIN/STM/exe_2nd ) );
    snl_invx05 \MAIN/STM/NS/U40  ( .ZN(\MAIN/STM/NS/n3341 ), .A(
        \MAIN/STM/NS/nst[1] ) );
    snl_ffqrnx1 \MAIN/STM/NS/est_reg[0]  ( .Q(\MAIN/STM/NS/nst[1] ), .D(
        \MAIN/STM/NS/nst[0] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nand03x0 \MAIN/STM/NS/U36  ( .ZN(\MAIN/STM/NS/n3343 ), .A(
        \MAIN/STM/NS/n3341 ), .B(\MAIN/STM/NS/n3338 ), .C(\MAIN/STM/NS/n3344 )
         );
    snl_invx05 \MAIN/STM/NS/U37  ( .ZN(\MAIN/STM/NS/n3340 ), .A(
        \MAIN/STM/exe_1st ) );
    snl_nand02x1 \MAIN/STM/NS/U39  ( .ZN(\MAIN/STM/NS/n3342 ), .A(st_exectl), 
        .B(\MAIN/reg_enable ) );
    snl_ffqrnx1 \MAIN/STM/NS/est_reg[1]  ( .Q(\MAIN/STM/NS/est[1] ), .D(
        \MAIN/STM/NS/nst[1] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \MAIN/STM/NS/U38  ( .ZN(\MAIN/STM/NS/n3338 ), .A(
        \MAIN/STM/NS/est[1] ) );
    snl_and02x1 \MAIN/STM/WS/U52  ( .Z(\MAIN/STM/WS/nwst[1] ), .A(
        \MAIN/STM/WS/ewst[0] ), .B(ph_lbend) );
    snl_nor02x1 \MAIN/STM/WS/U53  ( .ZN(\MAIN/STM/exec_eoc3 ), .A(
        \MAIN/STM/seq_doing ), .B(\MAIN/STM/WS/n3333 ) );
    snl_and02x1 \MAIN/STM/WS/U54  ( .Z(\MAIN/STM/exec_end3 ), .A(
        \MAIN/STM/WS/ewst[1] ), .B(\MAIN/STM/seq_doing ) );
    snl_nand12x1 \MAIN/STM/WS/U61  ( .ZN(\MAIN/STM/WS/n3336 ), .A(
        \MAIN/STM/WS/n3335 ), .B(\MAIN/STM/WS/n3333 ) );
    snl_ffqrnx1 \MAIN/STM/WS/ewst_reg[1]  ( .Q(\MAIN/STM/WS/ewst[1] ), .D(
        \MAIN/STM/WS/nwst[1] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \MAIN/STM/WS/U55  ( .ZN(\MAIN/STM/WS/n3333 ), .A(
        \MAIN/STM/WS/ewst[1] ) );
    snl_nor02x1 \MAIN/STM/WS/U56  ( .ZN(\MAIN/STM/WS/n3334 ), .A(
        \MAIN/STM/WS/ewst[0] ), .B(\MAIN/STM/WS/n3335 ) );
    snl_aoi022x1 \MAIN/STM/WS/U57  ( .ZN(\MAIN/STM/sa_start3 ), .A(
        \MAIN/STM/WS/n3334 ), .B(\MAIN/STM/WS/n3333 ), .C(
        \MAIN/STM/WS/ewst[0] ), .D(\MAIN/STM/WS/ewst[1] ) );
    snl_aoi113x0 \MAIN/STM/WS/U60  ( .ZN(\MAIN/STM/WS/n3335 ), .A(
        \MAIN/single_write ), .B(\MAIN/STM/WS/n3337 ), .C(st_exectl), .D(
        \MAIN/STM/exe_1st_w ), .E(\MAIN/STM/exe_2nd_w ) );
    snl_muxi21x1 \MAIN/STM/WS/U58  ( .ZN(phlbdir), .A(\MAIN/STM/WS/n3336 ), 
        .B(ph_lbend), .S(\MAIN/STM/WS/ewst[0] ) );
    snl_invx05 \MAIN/STM/WS/U59  ( .ZN(\MAIN/STM/WS/n3337 ), .A(
        \MAIN/seq_enable ) );
    snl_ffqrnx1 \MAIN/STM/WS/ewst_reg[0]  ( .Q(\MAIN/STM/WS/ewst[0] ), .D(
        phlbdir), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_ffqrnx1 \MAIN/STM/WS/exe_err_reg  ( .Q(\MAIN/STM/exe_err3 ), .D(
        ph_lberr), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nand13x1 \MAIN/STM/RS/U52  ( .ZN(\MAIN/STM/sa_start2 ), .A(
        \MAIN/STM/exec_eoc2 ), .B(\MAIN/STM/RS/n3324 ), .C(\MAIN/STM/RS/n3325 
        ) );
    snl_oai012x1 \MAIN/STM/RS/U53  ( .ZN(\MAIN/STM/RS/nrst[0] ), .A(
        \MAIN/STM/RS/n3326 ), .B(\MAIN/STM/RS/n3327 ), .C(\MAIN/STM/RS/n3328 )
         );
    snl_aoi012x1 \MAIN/STM/RS/U54  ( .ZN(\MAIN/STM/RS/n3326 ), .A(
        \MAIN/STM/RS/n3324 ), .B(\MAIN/STM/RS/n3329 ), .C(\MAIN/STM/exec_end2 
        ) );
    snl_nor02x1 \MAIN/STM/RS/U61  ( .ZN(\MAIN/STM/exec_eoc2 ), .A(
        \MAIN/STM/RS/n3329 ), .B(\MAIN/STM/seq_doing ) );
    snl_ffqrnx1 \MAIN/STM/RS/erst_reg[0]  ( .Q(\MAIN/STM/RS/erst[0] ), .D(
        \MAIN/STM/RS/nrst[0] ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_invx05 \MAIN/STM/RS/U55  ( .ZN(\MAIN/STM/RS/n3329 ), .A(
        \MAIN/STM/RS/erst[1] ) );
    snl_ffqrnx1 \MAIN/STM/RS/exe_error_reg  ( .Q(\MAIN/STM/exe_err2 ), .D(
        ph_lberr), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nand02x1 \MAIN/STM/RS/U56  ( .ZN(\MAIN/STM/RS/n3330 ), .A(st_exectl), 
        .B(\MAIN/single_read ) );
    snl_invx05 \MAIN/STM/RS/U57  ( .ZN(\MAIN/STM/RS/n3324 ), .A(
        \MAIN/STM/RS/erst[0] ) );
    snl_nor03x0 \MAIN/STM/RS/U60  ( .ZN(\MAIN/STM/RS/n3332 ), .A(
        \MAIN/STM/RS/n3330 ), .B(\MAIN/STM/RS/erst[1] ), .C(\MAIN/seq_enable )
         );
    snl_invx05 \MAIN/STM/RS/U58  ( .ZN(\MAIN/STM/RS/n3331 ), .A(ph_lbend) );
    snl_invx05 \MAIN/STM/RS/U59  ( .ZN(\MAIN/STM/RS/n3327 ), .A(
        \MAIN/STM/exe_1st_r ) );
    snl_and02x1 \MAIN/STM/RS/U62  ( .Z(\MAIN/STM/exec_end2 ), .A(
        \MAIN/STM/seq_doing ), .B(\MAIN/STM/RS/erst[1] ) );
    snl_aoi022x1 \MAIN/STM/RS/U65  ( .ZN(\MAIN/STM/RS/n3328 ), .A(
        \MAIN/STM/RS/n3331 ), .B(\MAIN/STM/RS/erst[0] ), .C(
        \MAIN/STM/RS/n3332 ), .D(\MAIN/STM/RS/n3324 ) );
    snl_oai013x0 \MAIN/STM/RS/U64  ( .ZN(\MAIN/STM/RS/n3325 ), .A(
        \MAIN/STM/RS/n3330 ), .B(\MAIN/STM/RS/erst[1] ), .C(\MAIN/seq_enable ), 
        .D(\MAIN/STM/RS/n3327 ) );
    snl_ffqrnx1 \MAIN/STM/RS/erst_reg[1]  ( .Q(\MAIN/STM/RS/erst[1] ), .D(
        \MAIN/STM/bnolth ), .RN(\MAIN/n3611 ), .CP(SCLK) );
    snl_nor02x1 \MAIN/STM/RS/U63  ( .ZN(\MAIN/STM/bnolth ), .A(
        \MAIN/STM/RS/n3331 ), .B(\MAIN/STM/RS/n3324 ) );
    snl_invx05 \SAEXE/RFIO/phcont4_1/ph4dec_1/U7  ( .ZN(
        \SAEXE/RFIO/phcont4_1/ncnt[0] ), .A(\SAEXE/RFIO/phcont4_1/count[0] )
         );
    snl_aoi022x1 \SAEXE/RFIO/phcont4_1/ph4dec_1/U8  ( .ZN(
        \SAEXE/RFIO/phcont4_1/ncnt[1] ), .A(\SAEXE/RFIO/phcont4_1/count[0] ), 
        .B(\SAEXE/RFIO/phcont4_1/ph4dec_1/n14 ), .C(
        \SAEXE/RFIO/phcont4_1/ncnt[0] ), .D(\SAEXE/RFIO/phcont4_1/count[1] )
         );
    snl_invx05 \SAEXE/RFIO/phcont4_1/ph4dec_1/U9  ( .ZN(
        \SAEXE/RFIO/phcont4_1/ph4dec_1/n14 ), .A(
        \SAEXE/RFIO/phcont4_1/count[1] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add0/U7  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/c_last ), .A(
        \SADR/MAINSADR/addidxof/add0/n8600 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8601 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8602 ) );
    snl_nor05x1 \SADR/MAINSADR/addidxof/add0/U8  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/gp_out ), .A(
        \SADR/MAINSADR/addidxof/add0/n8603 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8600 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8604 ), .D(
        \SADR/MAINSADR/addidxof/add0/n8605 ), .E(
        \SADR/MAINSADR/addidxof/add0/n8606 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U13  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8616 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8615 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8617 ) );
    snl_and12x1 \SADR/MAINSADR/addidxof/add0/U14  ( .Z(
        \SADR/MAINSADR/addidxof/add0/n8618 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8603 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8619 ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add0/U21  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8619 ), .A(\SADR/MAINSADR/index[0] ), 
        .B(\SADR/MAINSADR/offset[0] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add0/U28  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8621 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8600 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add0/U33  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8614 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8617 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U34  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8603 ), .A(\SADR/MAINSADR/index[0] ), 
        .B(\SADR/MAINSADR/offset[0] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add0/U41  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8602 ), .A(\SADR/MAINSADR/index[4] ), 
        .B(\SADR/MAINSADR/offset[4] ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add0/U46  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8624 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8625 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8629 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add0/U26  ( .Z(
        \SADR/MAINSADR/addindoff[0] ), .A(1'b0), .B(
        \SADR/MAINSADR/addidxof/add0/n8618 ) );
    snl_ao01b2x0 \SADR/MAINSADR/addidxof/add0/U9  ( .Z(
        \SADR/MAINSADR/addidxof/gg_out[0] ), .A(
        \SADR/MAINSADR/addidxof/add0/n8606 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8607 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8608 ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add0/U12  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8612 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8613 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8614 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8615 ) );
    snl_oai013x0 \SADR/MAINSADR/addidxof/add0/U35  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8623 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8627 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8603 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8605 ), .D(
        \SADR/MAINSADR/addidxof/add0/n8628 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U27  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8600 ), .A(\SADR/MAINSADR/index[4] ), 
        .B(\SADR/MAINSADR/offset[4] ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add0/U40  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8601 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8623 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8630 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8611 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add0/U20  ( .Z(
        \SADR/MAINSADR/addindoff[1] ), .A(\SADR/MAINSADR/addidxof/add0/n8613 ), 
        .B(\SADR/MAINSADR/addidxof/add0/n8616 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U29  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8625 ), .A(\SADR/MAINSADR/index[2] ), 
        .B(\SADR/MAINSADR/offset[2] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add0/U47  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8620 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8628 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8604 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8631 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U10  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8609 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8608 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8606 ) );
    snl_aoi0b12x0 \SADR/MAINSADR/addidxof/add0/U15  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8607 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8620 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8621 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8602 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add0/U17  ( .Z(
        \SADR/MAINSADR/addindoff[4] ), .A(\SADR/MAINSADR/addidxof/add0/n8622 ), 
        .B(\SADR/MAINSADR/addidxof/add0/n8601 ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add0/U22  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8605 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8625 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8614 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U32  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8617 ), .A(\SADR/MAINSADR/index[1] ), 
        .B(\SADR/MAINSADR/offset[1] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add0/U39  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8611 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8631 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add0/U30  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8615 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8626 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U42  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8606 ), .A(\SADR/MAINSADR/index[5] ), 
        .B(\SADR/MAINSADR/offset[5] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add0/U45  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8613 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8603 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8627 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8619 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U11  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8610 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8611 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8604 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add0/U19  ( .Z(
        \SADR/MAINSADR/addindoff[2] ), .A(\SADR/MAINSADR/addidxof/add0/n8624 ), 
        .B(\SADR/MAINSADR/addidxof/add0/n8612 ) );
    snl_oa122x1 \SADR/MAINSADR/addidxof/add0/U25  ( .Z(
        \SADR/MAINSADR/addidxof/add0/n8628 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8619 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8605 ), .C(
        \SADR/MAINSADR/addidxof/add0/n8625 ), .D(
        \SADR/MAINSADR/addidxof/add0/n8626 ), .E(
        \SADR/MAINSADR/addidxof/add0/n8629 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add0/U37  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8630 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8604 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add0/U16  ( .Z(
        \SADR/MAINSADR/addindoff[5] ), .A(\SADR/MAINSADR/addidxof/add0/c_last 
        ), .B(\SADR/MAINSADR/addidxof/add0/n8609 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add0/U18  ( .Z(
        \SADR/MAINSADR/addindoff[3] ), .A(\SADR/MAINSADR/addidxof/add0/n8623 ), 
        .B(\SADR/MAINSADR/addidxof/add0/n8610 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add0/U36  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8604 ), .A(\SADR/MAINSADR/index[3] ), 
        .B(\SADR/MAINSADR/offset[3] ) );
    snl_and02x1 \SADR/MAINSADR/addidxof/add0/U43  ( .Z(
        \SADR/MAINSADR/addidxof/add0/n8608 ), .A(\SADR/MAINSADR/index[5] ), 
        .B(\SADR/MAINSADR/offset[5] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add0/U23  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8626 ), .A(\SADR/MAINSADR/index[1] ), 
        .B(\SADR/MAINSADR/offset[1] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add0/U24  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8627 ), .A(1'b0) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add0/U31  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8629 ), .A(\SADR/MAINSADR/index[2] ), 
        .B(\SADR/MAINSADR/offset[2] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add0/U38  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8631 ), .A(\SADR/MAINSADR/index[3] ), 
        .B(\SADR/MAINSADR/offset[3] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add0/U44  ( .ZN(
        \SADR/MAINSADR/addidxof/add0/n8622 ), .A(
        \SADR/MAINSADR/addidxof/add0/n8621 ), .B(
        \SADR/MAINSADR/addidxof/add0/n8602 ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add1/U7  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/c_last ), .A(
        \SADR/MAINSADR/addidxof/add1/n8568 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8569 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8570 ) );
    snl_nor05x1 \SADR/MAINSADR/addidxof/add1/U8  ( .ZN(
        \SADR/MAINSADR/addidxof/gp_out[1] ), .A(
        \SADR/MAINSADR/addidxof/add1/n8571 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8568 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8572 ), .D(
        \SADR/MAINSADR/addidxof/add1/n8573 ), .E(
        \SADR/MAINSADR/addidxof/add1/n8574 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U13  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8584 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8583 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8585 ) );
    snl_and12x1 \SADR/MAINSADR/addidxof/add1/U14  ( .Z(
        \SADR/MAINSADR/addidxof/add1/n8586 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8571 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8587 ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add1/U21  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8587 ), .A(\SADR/MAINSADR/index[6] ), 
        .B(\SADR/MAINSADR/offset[6] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add1/U28  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8589 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8568 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add1/U33  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8582 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8585 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U34  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8571 ), .A(\SADR/MAINSADR/index[6] ), 
        .B(\SADR/MAINSADR/offset[6] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add1/U41  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8570 ), .A(\SADR/MAINSADR/index[10] ), 
        .B(\SADR/MAINSADR/offset[10] ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add1/U46  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8592 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8593 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8597 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add1/U26  ( .Z(
        \SADR/MAINSADR/addindoff[6] ), .A(\SADR/MAINSADR/addidxof/gg_out[0] ), 
        .B(\SADR/MAINSADR/addidxof/add1/n8586 ) );
    snl_ao01b2x0 \SADR/MAINSADR/addidxof/add1/U9  ( .Z(
        \SADR/MAINSADR/addidxof/gg_out[1] ), .A(
        \SADR/MAINSADR/addidxof/add1/n8574 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8575 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8576 ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add1/U12  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8580 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8581 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8582 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8583 ) );
    snl_oai013x0 \SADR/MAINSADR/addidxof/add1/U35  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8591 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8595 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8571 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8573 ), .D(
        \SADR/MAINSADR/addidxof/add1/n8596 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U27  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8568 ), .A(\SADR/MAINSADR/index[10] ), 
        .B(\SADR/MAINSADR/offset[10] ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add1/U40  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8569 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8591 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8598 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8579 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add1/U20  ( .Z(
        \SADR/MAINSADR/addindoff[7] ), .A(\SADR/MAINSADR/addidxof/add1/n8581 ), 
        .B(\SADR/MAINSADR/addidxof/add1/n8584 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U29  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8593 ), .A(\SADR/MAINSADR/index[8] ), 
        .B(\SADR/MAINSADR/offset[8] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add1/U47  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8588 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8596 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8572 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8599 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U10  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8577 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8576 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8574 ) );
    snl_aoi0b12x0 \SADR/MAINSADR/addidxof/add1/U15  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8575 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8588 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8589 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8570 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add1/U17  ( .Z(
        \SADR/MAINSADR/addindoff[10] ), .A(\SADR/MAINSADR/addidxof/add1/n8590 
        ), .B(\SADR/MAINSADR/addidxof/add1/n8569 ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add1/U22  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8573 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8593 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8582 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U32  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8585 ), .A(\SADR/MAINSADR/index[7] ), 
        .B(\SADR/MAINSADR/offset[7] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add1/U39  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8579 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8599 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add1/U30  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8583 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8594 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U42  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8574 ), .A(\SADR/MAINSADR/index[11] ), 
        .B(\SADR/MAINSADR/offset[11] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add1/U45  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8581 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8571 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8595 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8587 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U11  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8578 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8579 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8572 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add1/U19  ( .Z(
        \SADR/MAINSADR/addindoff[8] ), .A(\SADR/MAINSADR/addidxof/add1/n8592 ), 
        .B(\SADR/MAINSADR/addidxof/add1/n8580 ) );
    snl_oa122x1 \SADR/MAINSADR/addidxof/add1/U25  ( .Z(
        \SADR/MAINSADR/addidxof/add1/n8596 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8587 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8573 ), .C(
        \SADR/MAINSADR/addidxof/add1/n8593 ), .D(
        \SADR/MAINSADR/addidxof/add1/n8594 ), .E(
        \SADR/MAINSADR/addidxof/add1/n8597 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add1/U37  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8598 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8572 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add1/U16  ( .Z(
        \SADR/MAINSADR/addindoff[11] ), .A(
        \SADR/MAINSADR/addidxof/add1/c_last ), .B(
        \SADR/MAINSADR/addidxof/add1/n8577 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add1/U18  ( .Z(
        \SADR/MAINSADR/addindoff[9] ), .A(\SADR/MAINSADR/addidxof/add1/n8591 ), 
        .B(\SADR/MAINSADR/addidxof/add1/n8578 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add1/U36  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8572 ), .A(\SADR/MAINSADR/index[9] ), 
        .B(\SADR/MAINSADR/offset[9] ) );
    snl_and02x1 \SADR/MAINSADR/addidxof/add1/U43  ( .Z(
        \SADR/MAINSADR/addidxof/add1/n8576 ), .A(\SADR/MAINSADR/index[11] ), 
        .B(\SADR/MAINSADR/offset[11] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add1/U23  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8594 ), .A(\SADR/MAINSADR/index[7] ), 
        .B(\SADR/MAINSADR/offset[7] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add1/U24  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8595 ), .A(
        \SADR/MAINSADR/addidxof/gg_out[0] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add1/U31  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8597 ), .A(\SADR/MAINSADR/index[8] ), 
        .B(\SADR/MAINSADR/offset[8] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add1/U38  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8599 ), .A(\SADR/MAINSADR/index[9] ), 
        .B(\SADR/MAINSADR/offset[9] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add1/U44  ( .ZN(
        \SADR/MAINSADR/addidxof/add1/n8590 ), .A(
        \SADR/MAINSADR/addidxof/add1/n8589 ), .B(
        \SADR/MAINSADR/addidxof/add1/n8570 ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add2/U7  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/c_last ), .A(
        \SADR/MAINSADR/addidxof/add2/n8536 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8537 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8538 ) );
    snl_nor05x1 \SADR/MAINSADR/addidxof/add2/U8  ( .ZN(
        \SADR/MAINSADR/addidxof/gp_out[2] ), .A(
        \SADR/MAINSADR/addidxof/add2/n8539 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8536 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8540 ), .D(
        \SADR/MAINSADR/addidxof/add2/n8541 ), .E(
        \SADR/MAINSADR/addidxof/add2/n8542 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U13  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8552 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8551 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8553 ) );
    snl_and12x1 \SADR/MAINSADR/addidxof/add2/U14  ( .Z(
        \SADR/MAINSADR/addidxof/add2/n8554 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8539 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8555 ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add2/U21  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8555 ), .A(\SADR/MAINSADR/index[12] ), 
        .B(\SADR/MAINSADR/offset[12] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add2/U28  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8557 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8536 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add2/U33  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8550 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8553 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U34  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8539 ), .A(\SADR/MAINSADR/index[12] ), 
        .B(\SADR/MAINSADR/offset[12] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add2/U41  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8538 ), .A(\SADR/MAINSADR/index[16] ), 
        .B(\SADR/MAINSADR/offset[16] ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add2/U46  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8560 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8561 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8565 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add2/U26  ( .Z(
        \SADR/MAINSADR/addindoff[12] ), .A(\SADR/MAINSADR/addidxof/cin_stg[1] 
        ), .B(\SADR/MAINSADR/addidxof/add2/n8554 ) );
    snl_ao01b2x0 \SADR/MAINSADR/addidxof/add2/U9  ( .Z(
        \SADR/MAINSADR/addidxof/gg_out[2] ), .A(
        \SADR/MAINSADR/addidxof/add2/n8542 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8543 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8544 ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add2/U12  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8548 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8549 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8550 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8551 ) );
    snl_oai013x0 \SADR/MAINSADR/addidxof/add2/U35  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8559 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8563 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8539 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8541 ), .D(
        \SADR/MAINSADR/addidxof/add2/n8564 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U27  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8536 ), .A(\SADR/MAINSADR/index[16] ), 
        .B(\SADR/MAINSADR/offset[16] ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add2/U40  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8537 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8559 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8566 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8547 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add2/U20  ( .Z(
        \SADR/MAINSADR/addindoff[13] ), .A(\SADR/MAINSADR/addidxof/add2/n8549 
        ), .B(\SADR/MAINSADR/addidxof/add2/n8552 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U29  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8561 ), .A(\SADR/MAINSADR/index[14] ), 
        .B(\SADR/MAINSADR/offset[14] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add2/U47  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8556 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8564 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8540 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8567 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U10  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8545 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8544 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8542 ) );
    snl_aoi0b12x0 \SADR/MAINSADR/addidxof/add2/U15  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8543 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8556 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8557 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8538 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add2/U17  ( .Z(
        \SADR/MAINSADR/addindoff[16] ), .A(\SADR/MAINSADR/addidxof/add2/n8558 
        ), .B(\SADR/MAINSADR/addidxof/add2/n8537 ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add2/U22  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8541 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8561 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8550 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U32  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8553 ), .A(\SADR/MAINSADR/index[13] ), 
        .B(\SADR/MAINSADR/offset[13] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add2/U39  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8547 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8567 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add2/U30  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8551 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8562 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U42  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8542 ), .A(\SADR/MAINSADR/index[17] ), 
        .B(\SADR/MAINSADR/offset[17] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add2/U45  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8549 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8539 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8563 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8555 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U11  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8546 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8547 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8540 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add2/U19  ( .Z(
        \SADR/MAINSADR/addindoff[14] ), .A(\SADR/MAINSADR/addidxof/add2/n8560 
        ), .B(\SADR/MAINSADR/addidxof/add2/n8548 ) );
    snl_oa122x1 \SADR/MAINSADR/addidxof/add2/U25  ( .Z(
        \SADR/MAINSADR/addidxof/add2/n8564 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8555 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8541 ), .C(
        \SADR/MAINSADR/addidxof/add2/n8561 ), .D(
        \SADR/MAINSADR/addidxof/add2/n8562 ), .E(
        \SADR/MAINSADR/addidxof/add2/n8565 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add2/U37  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8566 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8540 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add2/U16  ( .Z(
        \SADR/MAINSADR/addindoff[17] ), .A(
        \SADR/MAINSADR/addidxof/add2/c_last ), .B(
        \SADR/MAINSADR/addidxof/add2/n8545 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add2/U18  ( .Z(
        \SADR/MAINSADR/addindoff[15] ), .A(\SADR/MAINSADR/addidxof/add2/n8559 
        ), .B(\SADR/MAINSADR/addidxof/add2/n8546 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add2/U36  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8540 ), .A(\SADR/MAINSADR/index[15] ), 
        .B(\SADR/MAINSADR/offset[15] ) );
    snl_and02x1 \SADR/MAINSADR/addidxof/add2/U43  ( .Z(
        \SADR/MAINSADR/addidxof/add2/n8544 ), .A(\SADR/MAINSADR/index[17] ), 
        .B(\SADR/MAINSADR/offset[17] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add2/U23  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8562 ), .A(\SADR/MAINSADR/index[13] ), 
        .B(\SADR/MAINSADR/offset[13] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add2/U24  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8563 ), .A(
        \SADR/MAINSADR/addidxof/cin_stg[1] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add2/U31  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8565 ), .A(\SADR/MAINSADR/index[14] ), 
        .B(\SADR/MAINSADR/offset[14] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add2/U38  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8567 ), .A(\SADR/MAINSADR/index[15] ), 
        .B(\SADR/MAINSADR/offset[15] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add2/U44  ( .ZN(
        \SADR/MAINSADR/addidxof/add2/n8558 ), .A(
        \SADR/MAINSADR/addidxof/add2/n8557 ), .B(
        \SADR/MAINSADR/addidxof/add2/n8538 ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add3/U7  ( .ZN(
        \SADR/MAINSADR/addidxof/c_last ), .A(
        \SADR/MAINSADR/addidxof/add3/n8504 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8505 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8506 ) );
    snl_nor05x1 \SADR/MAINSADR/addidxof/add3/U8  ( .ZN(
        \SADR/MAINSADR/addidxof/gp_out[3] ), .A(
        \SADR/MAINSADR/addidxof/add3/n8507 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8504 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8508 ), .D(
        \SADR/MAINSADR/addidxof/add3/n8509 ), .E(
        \SADR/MAINSADR/addidxof/add3/n8510 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U13  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8520 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8519 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8521 ) );
    snl_and12x1 \SADR/MAINSADR/addidxof/add3/U14  ( .Z(
        \SADR/MAINSADR/addidxof/add3/n8522 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8507 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8523 ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add3/U21  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8523 ), .A(\SADR/MAINSADR/index[18] ), 
        .B(\SADR/MAINSADR/offset[18] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add3/U28  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8525 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8504 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add3/U33  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8518 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8521 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U34  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8507 ), .A(\SADR/MAINSADR/index[18] ), 
        .B(\SADR/MAINSADR/offset[18] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add3/U41  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8506 ), .A(\SADR/MAINSADR/index[22] ), 
        .B(\SADR/MAINSADR/offset[22] ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add3/U46  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8528 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8529 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8533 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add3/U26  ( .Z(
        \SADR/MAINSADR/addindoff[18] ), .A(\SADR/MAINSADR/addidxof/cin_stg[2] 
        ), .B(\SADR/MAINSADR/addidxof/add3/n8522 ) );
    snl_ao01b2x0 \SADR/MAINSADR/addidxof/add3/U9  ( .Z(
        \SADR/MAINSADR/addidxof/gg_out[3] ), .A(
        \SADR/MAINSADR/addidxof/add3/n8510 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8511 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8512 ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add3/U12  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8516 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8517 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8518 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8519 ) );
    snl_oai013x0 \SADR/MAINSADR/addidxof/add3/U35  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8527 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8531 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8507 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8509 ), .D(
        \SADR/MAINSADR/addidxof/add3/n8532 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U27  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8504 ), .A(\SADR/MAINSADR/index[22] ), 
        .B(\SADR/MAINSADR/offset[22] ) );
    snl_aoi012x1 \SADR/MAINSADR/addidxof/add3/U40  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8505 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8527 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8534 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8515 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add3/U20  ( .Z(
        \SADR/MAINSADR/addindoff[19] ), .A(\SADR/MAINSADR/addidxof/add3/n8517 
        ), .B(\SADR/MAINSADR/addidxof/add3/n8520 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U29  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8529 ), .A(\SADR/MAINSADR/index[20] ), 
        .B(\SADR/MAINSADR/offset[20] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add3/U47  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8524 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8532 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8508 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8535 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U10  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8513 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8512 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8510 ) );
    snl_aoi0b12x0 \SADR/MAINSADR/addidxof/add3/U15  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8511 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8524 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8525 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8506 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add3/U17  ( .Z(
        \SADR/MAINSADR/addindoff[22] ), .A(\SADR/MAINSADR/addidxof/add3/n8526 
        ), .B(\SADR/MAINSADR/addidxof/add3/n8505 ) );
    snl_nand12x1 \SADR/MAINSADR/addidxof/add3/U22  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8509 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8529 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8518 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U32  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8521 ), .A(\SADR/MAINSADR/index[19] ), 
        .B(\SADR/MAINSADR/offset[19] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add3/U39  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8515 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8535 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add3/U30  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8519 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8530 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U42  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8510 ), .A(\SADR/MAINSADR/index[23] ), 
        .B(\SADR/MAINSADR/offset[23] ) );
    snl_oai012x1 \SADR/MAINSADR/addidxof/add3/U45  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8517 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8507 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8531 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8523 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U11  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8514 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8515 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8508 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add3/U19  ( .Z(
        \SADR/MAINSADR/addindoff[20] ), .A(\SADR/MAINSADR/addidxof/add3/n8528 
        ), .B(\SADR/MAINSADR/addidxof/add3/n8516 ) );
    snl_oa122x1 \SADR/MAINSADR/addidxof/add3/U25  ( .Z(
        \SADR/MAINSADR/addidxof/add3/n8532 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8523 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8509 ), .C(
        \SADR/MAINSADR/addidxof/add3/n8529 ), .D(
        \SADR/MAINSADR/addidxof/add3/n8530 ), .E(
        \SADR/MAINSADR/addidxof/add3/n8533 ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add3/U37  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8534 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8508 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add3/U16  ( .Z(
        \SADR/MAINSADR/addindoff[23] ), .A(\SADR/MAINSADR/addidxof/c_last ), 
        .B(\SADR/MAINSADR/addidxof/add3/n8513 ) );
    snl_xor2x0 \SADR/MAINSADR/addidxof/add3/U18  ( .Z(
        \SADR/MAINSADR/addindoff[21] ), .A(\SADR/MAINSADR/addidxof/add3/n8527 
        ), .B(\SADR/MAINSADR/addidxof/add3/n8514 ) );
    snl_nor02x1 \SADR/MAINSADR/addidxof/add3/U36  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8508 ), .A(\SADR/MAINSADR/index[21] ), 
        .B(\SADR/MAINSADR/offset[21] ) );
    snl_and02x1 \SADR/MAINSADR/addidxof/add3/U43  ( .Z(
        \SADR/MAINSADR/addidxof/add3/n8512 ), .A(\SADR/MAINSADR/index[23] ), 
        .B(\SADR/MAINSADR/offset[23] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add3/U23  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8530 ), .A(\SADR/MAINSADR/index[19] ), 
        .B(\SADR/MAINSADR/offset[19] ) );
    snl_invx05 \SADR/MAINSADR/addidxof/add3/U24  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8531 ), .A(
        \SADR/MAINSADR/addidxof/cin_stg[2] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add3/U31  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8533 ), .A(\SADR/MAINSADR/index[20] ), 
        .B(\SADR/MAINSADR/offset[20] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add3/U38  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8535 ), .A(\SADR/MAINSADR/index[21] ), 
        .B(\SADR/MAINSADR/offset[21] ) );
    snl_nand02x1 \SADR/MAINSADR/addidxof/add3/U44  ( .ZN(
        \SADR/MAINSADR/addidxof/add3/n8526 ), .A(
        \SADR/MAINSADR/addidxof/add3/n8525 ), .B(
        \SADR/MAINSADR/addidxof/add3/n8506 ) );
    snl_and05x1 \SADR/MAINSADR/addsegoff/add0/U7  ( .Z(
        \SADR/MAINSADR/addsegoff/add0/gp_out ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8461 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8462 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8463 ), .D(
        \SADR/MAINSADR/addsegoff/add0/n8464 ), .E(
        \SADR/MAINSADR/addsegoff/add0/n8465 ) );
    snl_oai012x1 \SADR/MAINSADR/addsegoff/add0/U8  ( .ZN(
        \SADR/MAINSADR/addsegoff/gg_out[0] ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8466 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8467 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8468 ) );
    snl_and02x1 \SADR/MAINSADR/addsegoff/add0/U13  ( .Z(
        \SADR/MAINSADR/addsegoff/add0/n8481 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8482 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8461 ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/add0/U14  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8467 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8483 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8462 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8471 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U21  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8464 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8480 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8488 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U28  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8488 ), .A(\SADR/segbase[2] ), .B(
        \pgsdprlh[15] ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U33  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8494 ), .A(\SADR/segbase[0] ), .B(
        \pgsdprlh[13] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U34  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8461 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8494 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U41  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8496 ), .A(\SADR/segbase[4] ), .B(
        \pgsdprlh[17] ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U46  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8484 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8465 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8468 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U26  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8492 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8464 ) );
    snl_oai012x1 \SADR/MAINSADR/addsegoff/add0/U48  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8476 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8494 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8490 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8482 ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/add0/U9  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8469 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8470 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8462 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8471 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U12  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8479 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8478 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8480 ) );
    snl_oai013x0 \SADR/MAINSADR/addsegoff/add0/U35  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8486 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8490 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8494 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8492 ), .D(
        \SADR/MAINSADR/addsegoff/add0/n8491 ) );
    snl_or02x1 \SADR/MAINSADR/addsegoff/add0/U27  ( .Z(
        \SADR/MAINSADR/addsegoff/add0/n8462 ), .A(\SADR/segbase[4] ), .B(
        \pgsdprlh[17] ) );
    snl_ao012x1 \SADR/MAINSADR/addsegoff/add0/U40  ( .Z(
        \SADR/MAINSADR/addsegoff/add0/n8470 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8486 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8463 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8473 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U20  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8482 ), .A(\SADR/segbase[0] ), .B(
        \pgsdprlh[13] ) );
    snl_nand12x1 \SADR/MAINSADR/addsegoff/add0/U49  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8487 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8488 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8493 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U29  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8478 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8489 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U47  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8485 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8462 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8496 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U10  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8472 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8473 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8474 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add0/U15  ( .Z(\SADR/sadr[15] ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8484 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8469 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add0/U17  ( .Z(\SADR/sadr[13] ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8486 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8472 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U22  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8489 ), .A(\SADR/segbase[1] ), .B(
        \pgsdprlh[14] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U32  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8477 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8480 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U39  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8473 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8495 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U30  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8493 ), .A(\SADR/segbase[2] ), .B(
        \pgsdprlh[15] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U42  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8471 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8496 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U45  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8468 ), .A(\SADR/segbase[5] ), .B(
        \pgsdprlh[18] ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/add0/U11  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8475 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8476 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8477 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8478 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add0/U19  ( .Z(\SADR/sadr[11] ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8476 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8479 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add0/U25  ( .Z(\SADR/sadr[10] ), .A(
        1'b0), .B(\SADR/MAINSADR/addsegoff/add0/n8481 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U37  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8463 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8474 ) );
    snl_oai012x1 \SADR/MAINSADR/addsegoff/add0/U50  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8483 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8491 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8474 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8495 ) );
    snl_xnor2x0 \SADR/MAINSADR/addsegoff/add0/U16  ( .ZN(\SADR/sadr[14] ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8485 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8470 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add0/U18  ( .Z(\SADR/sadr[12] ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8487 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8475 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U36  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8474 ), .A(\SADR/segbase[3] ), .B(
        \pgsdprlh[16] ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U43  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8466 ), .A(\SADR/segbase[5] ), .B(
        \pgsdprlh[18] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U23  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8490 ), .A(1'b0) );
    snl_oa122x1 \SADR/MAINSADR/addsegoff/add0/U24  ( .Z(
        \SADR/MAINSADR/addsegoff/add0/n8491 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8482 ), .B(
        \SADR/MAINSADR/addsegoff/add0/n8492 ), .C(
        \SADR/MAINSADR/addsegoff/add0/n8488 ), .D(
        \SADR/MAINSADR/addsegoff/add0/n8489 ), .E(
        \SADR/MAINSADR/addsegoff/add0/n8493 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add0/U31  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8480 ), .A(\SADR/segbase[1] ), .B(
        \pgsdprlh[14] ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add0/U38  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8495 ), .A(\SADR/segbase[3] ), .B(
        \pgsdprlh[16] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add0/U44  ( .ZN(
        \SADR/MAINSADR/addsegoff/add0/n8465 ), .A(
        \SADR/MAINSADR/addsegoff/add0/n8466 ) );
    snl_and05x1 \SADR/MAINSADR/addsegoff/add1/U7  ( .Z(
        \SADR/MAINSADR/addsegoff/gp_out[1] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8425 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8426 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8427 ), .D(
        \SADR/MAINSADR/addsegoff/add1/n8428 ), .E(
        \SADR/MAINSADR/addsegoff/add1/n8429 ) );
    snl_oai012x1 \SADR/MAINSADR/addsegoff/add1/U8  ( .ZN(
        \SADR/MAINSADR/addsegoff/gg_out[1] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8430 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8431 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8432 ) );
    snl_and02x1 \SADR/MAINSADR/addsegoff/add1/U13  ( .Z(
        \SADR/MAINSADR/addsegoff/add1/n8445 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8446 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8425 ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/add1/U14  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8431 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8447 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8426 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8435 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U21  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8428 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8444 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8452 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U28  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8452 ), .A(\SADR/segbase[8] ), .B(
        \pgsdprlh[21] ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U33  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8458 ), .A(\SADR/segbase[6] ), .B(
        \pgsdprlh[19] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U34  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8425 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8458 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U41  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8460 ), .A(\SADR/segbase[10] ), .B(
        \pgsdprlh[23] ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U46  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8448 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8429 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8432 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U26  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8456 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8428 ) );
    snl_oai012x1 \SADR/MAINSADR/addsegoff/add1/U48  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8440 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8458 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8454 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8446 ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/add1/U9  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8433 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8434 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8426 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8435 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U12  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8443 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8442 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8444 ) );
    snl_oai013x0 \SADR/MAINSADR/addsegoff/add1/U35  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8450 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8454 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8458 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8456 ), .D(
        \SADR/MAINSADR/addsegoff/add1/n8455 ) );
    snl_or02x1 \SADR/MAINSADR/addsegoff/add1/U27  ( .Z(
        \SADR/MAINSADR/addsegoff/add1/n8426 ), .A(\SADR/segbase[10] ), .B(
        \pgsdprlh[23] ) );
    snl_ao012x1 \SADR/MAINSADR/addsegoff/add1/U40  ( .Z(
        \SADR/MAINSADR/addsegoff/add1/n8434 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8450 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8427 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8437 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U20  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8446 ), .A(\SADR/segbase[6] ), .B(
        \pgsdprlh[19] ) );
    snl_nand12x1 \SADR/MAINSADR/addsegoff/add1/U49  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8451 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8452 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8457 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U29  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8442 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8453 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U47  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8449 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8426 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8460 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U10  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8436 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8437 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8438 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add1/U15  ( .Z(\SADR/sadr[21] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8448 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8433 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add1/U17  ( .Z(\SADR/sadr[19] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8450 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8436 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U22  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8453 ), .A(\SADR/segbase[7] ), .B(
        \pgsdprlh[20] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U32  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8441 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8444 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U39  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8437 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8459 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U30  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8457 ), .A(\SADR/segbase[8] ), .B(
        \pgsdprlh[21] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U42  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8435 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8460 ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U45  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8432 ), .A(\SADR/segbase[11] ), .B(1'b0
        ) );
    snl_aoi012x1 \SADR/MAINSADR/addsegoff/add1/U11  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8439 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8440 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8441 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8442 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add1/U19  ( .Z(\SADR/sadr[17] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8440 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8443 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add1/U25  ( .Z(\SADR/sadr[16] ), .A(
        \SADR/MAINSADR/addsegoff/gg_out[0] ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8445 ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U37  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8427 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8438 ) );
    snl_oai012x1 \SADR/MAINSADR/addsegoff/add1/U50  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8447 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8455 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8438 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8459 ) );
    snl_xnor2x0 \SADR/MAINSADR/addsegoff/add1/U16  ( .ZN(\SADR/sadr[20] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8449 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8434 ) );
    snl_xor2x0 \SADR/MAINSADR/addsegoff/add1/U18  ( .Z(\SADR/sadr[18] ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8451 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8439 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U36  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8438 ), .A(\SADR/segbase[9] ), .B(
        \pgsdprlh[22] ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U43  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8430 ), .A(\SADR/segbase[11] ), .B(1'b0
        ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U23  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8454 ), .A(
        \SADR/MAINSADR/addsegoff/gg_out[0] ) );
    snl_oa122x1 \SADR/MAINSADR/addsegoff/add1/U24  ( .Z(
        \SADR/MAINSADR/addsegoff/add1/n8455 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8446 ), .B(
        \SADR/MAINSADR/addsegoff/add1/n8456 ), .C(
        \SADR/MAINSADR/addsegoff/add1/n8452 ), .D(
        \SADR/MAINSADR/addsegoff/add1/n8453 ), .E(
        \SADR/MAINSADR/addsegoff/add1/n8457 ) );
    snl_nor02x1 \SADR/MAINSADR/addsegoff/add1/U31  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8444 ), .A(\SADR/segbase[7] ), .B(
        \pgsdprlh[20] ) );
    snl_nand02x1 \SADR/MAINSADR/addsegoff/add1/U38  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8459 ), .A(\SADR/segbase[9] ), .B(
        \pgsdprlh[22] ) );
    snl_invx05 \SADR/MAINSADR/addsegoff/add1/U44  ( .ZN(
        \SADR/MAINSADR/addsegoff/add1/n8429 ), .A(
        \SADR/MAINSADR/addsegoff/add1/n8430 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc1/inc4_1/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/gp_out[0] ), .A(\SADR/MAINSADR/oddadd[3] ), .B(
        \SADR/MAINSADR/oddadd[0] ), .C(\SADR/MAINSADR/oddadd[1] ), .D(
        \SADR/MAINSADR/oddadd[2] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_1/U8  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_1/n8422 ), .A(\SADR/MAINSADR/oddadd[0] ), 
        .B(1'b1) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_1/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p1[0] ), .A(\SADR/MAINSADR/oddadd[0] ), .B(1'b1)
         );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_1/U14  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_1/n8424 ), .A(\SADR/MAINSADR/oddadd[2] ), 
        .B(\SADR/MAINSADR/adrinc1/inc4_1/n8423 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc1/inc4_1/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_1/n8423 ), .A(
        \SADR/MAINSADR/adrinc1/inc4_1/n8422 ), .B(\SADR/MAINSADR/oddadd[1] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_1/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[1] ), .A(\SADR/MAINSADR/oddadd[1] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_1/n8422 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_1/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[3] ), .A(\SADR/MAINSADR/oddadd[3] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_1/n8424 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_1/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p1[2] ), .A(\SADR/MAINSADR/oddadd[2] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_1/n8423 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc1/inc4_6/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_6/gp_out ), .A(\SADR/MAINSADR/oddadd[23] ), 
        .B(\SADR/MAINSADR/oddadd[20] ), .C(\SADR/MAINSADR/oddadd[21] ), .D(
        \SADR/MAINSADR/oddadd[22] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_6/U8  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_6/n8419 ), .A(\SADR/MAINSADR/oddadd[20] ), 
        .B(\SADR/MAINSADR/adrinc1/gg_out[4] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_6/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p1[20] ), .A(\SADR/MAINSADR/oddadd[20] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[4] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_6/U14  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_6/n8421 ), .A(\SADR/MAINSADR/oddadd[22] ), 
        .B(\SADR/MAINSADR/adrinc1/inc4_6/n8420 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc1/inc4_6/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_6/n8420 ), .A(
        \SADR/MAINSADR/adrinc1/inc4_6/n8419 ), .B(\SADR/MAINSADR/oddadd[21] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_6/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[21] ), .A(\SADR/MAINSADR/oddadd[21] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_6/n8419 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_6/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[23] ), .A(\SADR/MAINSADR/oddadd[23] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_6/n8421 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_6/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p1[22] ), .A(\SADR/MAINSADR/oddadd[22] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_6/n8420 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc1/inc4_2/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/gp_out[1] ), .A(\SADR/MAINSADR/oddadd[7] ), .B(
        \SADR/MAINSADR/oddadd[4] ), .C(\SADR/MAINSADR/oddadd[5] ), .D(
        \SADR/MAINSADR/oddadd[6] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_2/U8  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_2/n8416 ), .A(\SADR/MAINSADR/oddadd[4] ), 
        .B(\SADR/MAINSADR/adrinc1/gp_out[0] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_2/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p1[4] ), .A(\SADR/MAINSADR/oddadd[4] ), .B(
        \SADR/MAINSADR/adrinc1/gp_out[0] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_2/U14  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_2/n8418 ), .A(\SADR/MAINSADR/oddadd[6] ), 
        .B(\SADR/MAINSADR/adrinc1/inc4_2/n8417 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc1/inc4_2/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_2/n8417 ), .A(
        \SADR/MAINSADR/adrinc1/inc4_2/n8416 ), .B(\SADR/MAINSADR/oddadd[5] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_2/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[5] ), .A(\SADR/MAINSADR/oddadd[5] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_2/n8416 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_2/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[7] ), .A(\SADR/MAINSADR/oddadd[7] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_2/n8418 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_2/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p1[6] ), .A(\SADR/MAINSADR/oddadd[6] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_2/n8417 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc1/inc4_3/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/gp_out[2] ), .A(\SADR/MAINSADR/oddadd[11] ), 
        .B(\SADR/MAINSADR/oddadd[8] ), .C(\SADR/MAINSADR/oddadd[9] ), .D(
        \SADR/MAINSADR/oddadd[10] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_3/U8  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_3/n8413 ), .A(\SADR/MAINSADR/oddadd[8] ), 
        .B(\SADR/MAINSADR/adrinc1/gg_out[1] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_3/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p1[8] ), .A(\SADR/MAINSADR/oddadd[8] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[1] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_3/U14  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_3/n8415 ), .A(\SADR/MAINSADR/oddadd[10] ), 
        .B(\SADR/MAINSADR/adrinc1/inc4_3/n8414 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc1/inc4_3/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_3/n8414 ), .A(
        \SADR/MAINSADR/adrinc1/inc4_3/n8413 ), .B(\SADR/MAINSADR/oddadd[9] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_3/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[9] ), .A(\SADR/MAINSADR/oddadd[9] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_3/n8413 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_3/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[11] ), .A(\SADR/MAINSADR/oddadd[11] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_3/n8415 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_3/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p1[10] ), .A(\SADR/MAINSADR/oddadd[10] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_3/n8414 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc1/inc4_4/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/gp_out[3] ), .A(\SADR/MAINSADR/oddadd[15] ), 
        .B(\SADR/MAINSADR/oddadd[12] ), .C(\SADR/MAINSADR/oddadd[13] ), .D(
        \SADR/MAINSADR/oddadd[14] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_4/U8  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_4/n8410 ), .A(\SADR/MAINSADR/oddadd[12] ), 
        .B(\SADR/MAINSADR/adrinc1/gg_out[2] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_4/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p1[12] ), .A(\SADR/MAINSADR/oddadd[12] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[2] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_4/U14  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_4/n8412 ), .A(\SADR/MAINSADR/oddadd[14] ), 
        .B(\SADR/MAINSADR/adrinc1/inc4_4/n8411 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc1/inc4_4/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_4/n8411 ), .A(
        \SADR/MAINSADR/adrinc1/inc4_4/n8410 ), .B(\SADR/MAINSADR/oddadd[13] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_4/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[13] ), .A(\SADR/MAINSADR/oddadd[13] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_4/n8410 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_4/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[15] ), .A(\SADR/MAINSADR/oddadd[15] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_4/n8412 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_4/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p1[14] ), .A(\SADR/MAINSADR/oddadd[14] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_4/n8411 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc1/inc4_5/U7  ( .Z(
        \SADR/MAINSADR/adrinc1/gp_out[4] ), .A(\SADR/MAINSADR/oddadd[19] ), 
        .B(\SADR/MAINSADR/oddadd[16] ), .C(\SADR/MAINSADR/oddadd[17] ), .D(
        \SADR/MAINSADR/oddadd[18] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_5/U8  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_5/n8407 ), .A(\SADR/MAINSADR/oddadd[16] ), 
        .B(\SADR/MAINSADR/adrinc1/gg_out[3] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_5/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p1[16] ), .A(\SADR/MAINSADR/oddadd[16] ), .B(
        \SADR/MAINSADR/adrinc1/gg_out[3] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc1/inc4_5/U14  ( .ZN(
        \SADR/MAINSADR/adrinc1/inc4_5/n8409 ), .A(\SADR/MAINSADR/oddadd[18] ), 
        .B(\SADR/MAINSADR/adrinc1/inc4_5/n8408 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc1/inc4_5/U9  ( .Z(
        \SADR/MAINSADR/adrinc1/inc4_5/n8408 ), .A(
        \SADR/MAINSADR/adrinc1/inc4_5/n8407 ), .B(\SADR/MAINSADR/oddadd[17] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_5/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[17] ), .A(\SADR/MAINSADR/oddadd[17] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_5/n8407 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc1/inc4_5/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p1[19] ), .A(\SADR/MAINSADR/oddadd[19] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_5/n8409 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc1/inc4_5/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p1[18] ), .A(\SADR/MAINSADR/oddadd[18] ), .B(
        \SADR/MAINSADR/adrinc1/inc4_5/n8408 ) );
    snl_oai022x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U10  ( .ZN(
        \SADR/MAINSADR/adrcmp1/ggfl[3] ), .A(\pgsdprlh[23] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8390 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8391 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8392 ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U12  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8395 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8396 ), .B(\pgsdprlh[22] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U13  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8391 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8390 ), .B(\pgsdprlh[23] ) );
    snl_nor04x0 \SADR/MAINSADR/adrcmp1/cmp4_3/U14  ( .ZN(
        \SADR/MAINSADR/adrcmp1/geq[3] ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8397 ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8398 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8399 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8400 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_3/U21  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8402 ), .A(\pgsdprlh[20] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_3/U15  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8401 ), .A(\SADR/lmtaddr[13] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_3/U20  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8392 ), .A(\SADR/lmtaddr[15] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U17  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8396 ), .A(\pgsdprlh[21] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8394 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8393 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8401 ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_3/U22  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8397 ), .A(\SADR/lmtaddr[14] ), .B(
        \pgsdprlh[22] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U11  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8393 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8394 ), .B(\pgsdprlh[21] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U19  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8390 ), .A(\pgsdprlh[22] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8396 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8395 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8403 ) );
    snl_oai012x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U25  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8398 ), .A(\SADR/lmtaddr[12] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8402 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8394 ) );
    snl_nand02x1 \SADR/MAINSADR/adrcmp1/cmp4_3/U16  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8394 ), .A(\SADR/lmtaddr[12] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8402 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_3/U18  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8403 ), .A(\SADR/lmtaddr[14] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_3/U23  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8399 ), .A(\SADR/lmtaddr[13] ), .B(
        \pgsdprlh[21] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_3/U24  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_3/n8400 ), .A(\SADR/lmtaddr[15] ), .B(
        \pgsdprlh[23] ) );
    snl_oai022x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U10  ( .ZN(
        \SADR/MAINSADR/adrcmp1/ggfl[1] ), .A(\pgsdprlh[15] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8376 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8377 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8378 ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U12  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8381 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8382 ), .B(\pgsdprlh[14] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U13  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8377 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8376 ), .B(\pgsdprlh[15] ) );
    snl_nor04x0 \SADR/MAINSADR/adrcmp1/cmp4_1/U14  ( .ZN(
        \SADR/MAINSADR/adrcmp1/geq[1] ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8383 ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8384 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8385 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8386 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_1/U21  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8388 ), .A(\pgsdprlh[12] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_1/U15  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8387 ), .A(\SADR/lmtaddr[5] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_1/U20  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8378 ), .A(\SADR/lmtaddr[7] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U17  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8382 ), .A(\pgsdprlh[13] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8380 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8379 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8387 ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_1/U22  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8383 ), .A(\SADR/lmtaddr[6] ), .B(
        \pgsdprlh[14] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U11  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8379 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8380 ), .B(\pgsdprlh[13] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U19  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8376 ), .A(\pgsdprlh[14] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8382 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8381 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8389 ) );
    snl_oai012x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U25  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8384 ), .A(\SADR/lmtaddr[4] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8388 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8380 ) );
    snl_nand02x1 \SADR/MAINSADR/adrcmp1/cmp4_1/U16  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8380 ), .A(\SADR/lmtaddr[4] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8388 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_1/U18  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8389 ), .A(\SADR/lmtaddr[6] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_1/U23  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8385 ), .A(\SADR/lmtaddr[5] ), .B(
        \pgsdprlh[13] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_1/U24  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_1/n8386 ), .A(\SADR/lmtaddr[7] ), .B(
        \pgsdprlh[15] ) );
    snl_oai022x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U10  ( .ZN(
        \SADR/MAINSADR/adrcmp1/ggfl[0] ), .A(\pgsdprlh[11] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8362 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8363 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8364 ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U12  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8367 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8368 ), .B(\pgsdprlh[10] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U13  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8363 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8362 ), .B(\pgsdprlh[11] ) );
    snl_nor04x0 \SADR/MAINSADR/adrcmp1/cmp4_0/U14  ( .ZN(
        \SADR/MAINSADR/adrcmp1/geq[0] ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8369 ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8370 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8371 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8372 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_0/U21  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8374 ), .A(\pgsdprlh[8] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_0/U15  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8373 ), .A(\SADR/lmtaddr[1] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_0/U20  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8364 ), .A(\SADR/lmtaddr[3] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U17  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8368 ), .A(\pgsdprlh[9] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8366 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8365 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8373 ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_0/U22  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8369 ), .A(\SADR/lmtaddr[2] ), .B(
        \pgsdprlh[10] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U11  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8365 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8366 ), .B(\pgsdprlh[9] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U19  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8362 ), .A(\pgsdprlh[10] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8368 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8367 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8375 ) );
    snl_oai012x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U25  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8370 ), .A(\SADR/lmtaddr[0] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8374 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8366 ) );
    snl_nand02x1 \SADR/MAINSADR/adrcmp1/cmp4_0/U16  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8366 ), .A(\SADR/lmtaddr[0] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8374 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_0/U18  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8375 ), .A(\SADR/lmtaddr[2] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_0/U23  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8371 ), .A(\SADR/lmtaddr[1] ), .B(
        \pgsdprlh[9] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_0/U24  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_0/n8372 ), .A(\SADR/lmtaddr[3] ), .B(
        \pgsdprlh[11] ) );
    snl_oai022x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U10  ( .ZN(
        \SADR/MAINSADR/adrcmp1/ggfl[2] ), .A(\pgsdprlh[19] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8348 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8349 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8350 ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U12  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8353 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8354 ), .B(\pgsdprlh[18] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U13  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8349 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8348 ), .B(\pgsdprlh[19] ) );
    snl_nor04x0 \SADR/MAINSADR/adrcmp1/cmp4_2/U14  ( .ZN(
        \SADR/MAINSADR/adrcmp1/geq[2] ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8355 ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8356 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8357 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8358 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_2/U21  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8360 ), .A(\pgsdprlh[16] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_2/U15  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8359 ), .A(\SADR/lmtaddr[9] ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_2/U20  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8350 ), .A(\SADR/lmtaddr[11] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U17  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8354 ), .A(\pgsdprlh[17] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8352 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8351 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8359 ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_2/U22  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8355 ), .A(\SADR/lmtaddr[10] ), .B(
        \pgsdprlh[18] ) );
    snl_and02x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U11  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8351 ), .A(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8352 ), .B(\pgsdprlh[17] ) );
    snl_oa022x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U19  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8348 ), .A(\pgsdprlh[18] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8354 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8353 ), .D(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8361 ) );
    snl_oai012x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U25  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8356 ), .A(\SADR/lmtaddr[8] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8360 ), .C(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8352 ) );
    snl_nand02x1 \SADR/MAINSADR/adrcmp1/cmp4_2/U16  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8352 ), .A(\SADR/lmtaddr[8] ), .B(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8360 ) );
    snl_invx05 \SADR/MAINSADR/adrcmp1/cmp4_2/U18  ( .ZN(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8361 ), .A(\SADR/lmtaddr[10] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_2/U23  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8357 ), .A(\SADR/lmtaddr[9] ), .B(
        \pgsdprlh[17] ) );
    snl_xor2x0 \SADR/MAINSADR/adrcmp1/cmp4_2/U24  ( .Z(
        \SADR/MAINSADR/adrcmp1/cmp4_2/n8358 ), .A(\SADR/lmtaddr[11] ), .B(
        \pgsdprlh[19] ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec1/dec4_1/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m1[0] ), .A(\SADR/MAINSADR/oddadd[0] ), .B(1'b0), 
        .C(\SADR/MAINSADR/adrdec1/dec4_1/n8342 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec1/dec4_1/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/gg_out[0] ), .A(\SADR/MAINSADR/oddadd[0] ), .B(
        \SADR/MAINSADR/oddadd[3] ), .C(\SADR/MAINSADR/oddadd[1] ), .D(
        \SADR/MAINSADR/oddadd[2] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec1/dec4_1/U13  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_1/n8346 ), .A(
        \SADR/MAINSADR/adrdec1/dec4_1/n8342 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_1/n8345 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_1/U14  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_1/n8344 ), .A(\SADR/MAINSADR/oddadd[3] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec1/dec4_1/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[3] ), .A(1'b0), .B(
        \SADR/MAINSADR/adrdec1/gg_out[0] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_1/n8343 ), .D(
        \SADR/MAINSADR/adrdec1/dec4_1/n8344 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_1/U12  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_1/n8342 ), .A(1'b0), .B(
        \SADR/MAINSADR/oddadd[0] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec1/dec4_1/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[1] ), .A(\SADR/MAINSADR/adrdec1/dec4_1/n8342 
        ), .B(\SADR/MAINSADR/adrdec1/dec4_1/n8345 ), .C(
        \SADR/MAINSADR/adrdec1/dec4_1/n8346 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_1/U15  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_1/n8345 ), .A(\SADR/MAINSADR/oddadd[1] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_1/U11  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_1/n8343 ), .A(\SADR/MAINSADR/oddadd[2] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_1/n8346 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec1/dec4_1/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[2] ), .A(\SADR/MAINSADR/oddadd[2] ), .B(
        \SADR/MAINSADR/adrdec1/dec4_1/n8346 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec1/dec4_2/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m1[4] ), .A(\SADR/MAINSADR/oddadd[4] ), .B(
        \SADR/MAINSADR/adrdec1/gg_out[0] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_2/n8337 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec1/dec4_2/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/gg_out[1] ), .A(\SADR/MAINSADR/oddadd[4] ), .B(
        \SADR/MAINSADR/oddadd[7] ), .C(\SADR/MAINSADR/oddadd[5] ), .D(
        \SADR/MAINSADR/oddadd[6] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec1/dec4_2/U13  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_2/n8341 ), .A(
        \SADR/MAINSADR/adrdec1/dec4_2/n8337 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_2/n8340 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_2/U14  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_2/n8339 ), .A(\SADR/MAINSADR/oddadd[7] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec1/dec4_2/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[7] ), .A(\SADR/MAINSADR/adrdec1/gg_out[0] ), 
        .B(\SADR/MAINSADR/adrdec1/gg_out[1] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_2/n8338 ), .D(
        \SADR/MAINSADR/adrdec1/dec4_2/n8339 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_2/U12  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_2/n8337 ), .A(
        \SADR/MAINSADR/adrdec1/gg_out[0] ), .B(\SADR/MAINSADR/oddadd[4] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec1/dec4_2/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[5] ), .A(\SADR/MAINSADR/adrdec1/dec4_2/n8337 
        ), .B(\SADR/MAINSADR/adrdec1/dec4_2/n8340 ), .C(
        \SADR/MAINSADR/adrdec1/dec4_2/n8341 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_2/U15  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_2/n8340 ), .A(\SADR/MAINSADR/oddadd[5] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_2/U11  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_2/n8338 ), .A(\SADR/MAINSADR/oddadd[6] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_2/n8341 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec1/dec4_2/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[6] ), .A(\SADR/MAINSADR/oddadd[6] ), .B(
        \SADR/MAINSADR/adrdec1/dec4_2/n8341 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec1/dec4_3/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m1[8] ), .A(\SADR/MAINSADR/oddadd[8] ), .B(
        \SADR/MAINSADR/adrdec1/gcarry[1] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_3/n8332 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec1/dec4_3/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/gg_out[2] ), .A(\SADR/MAINSADR/oddadd[8] ), .B(
        \SADR/MAINSADR/oddadd[11] ), .C(\SADR/MAINSADR/oddadd[9] ), .D(
        \SADR/MAINSADR/oddadd[10] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec1/dec4_3/U13  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_3/n8336 ), .A(
        \SADR/MAINSADR/adrdec1/dec4_3/n8332 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_3/n8335 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_3/U14  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_3/n8334 ), .A(\SADR/MAINSADR/oddadd[11] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec1/dec4_3/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[11] ), .A(\SADR/MAINSADR/adrdec1/gcarry[1] ), 
        .B(\SADR/MAINSADR/adrdec1/gg_out[2] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_3/n8333 ), .D(
        \SADR/MAINSADR/adrdec1/dec4_3/n8334 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_3/U12  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_3/n8332 ), .A(
        \SADR/MAINSADR/adrdec1/gcarry[1] ), .B(\SADR/MAINSADR/oddadd[8] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec1/dec4_3/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[9] ), .A(\SADR/MAINSADR/adrdec1/dec4_3/n8332 
        ), .B(\SADR/MAINSADR/adrdec1/dec4_3/n8335 ), .C(
        \SADR/MAINSADR/adrdec1/dec4_3/n8336 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_3/U15  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_3/n8335 ), .A(\SADR/MAINSADR/oddadd[9] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_3/U11  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_3/n8333 ), .A(\SADR/MAINSADR/oddadd[10] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_3/n8336 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec1/dec4_3/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[10] ), .A(\SADR/MAINSADR/oddadd[10] ), .B(
        \SADR/MAINSADR/adrdec1/dec4_3/n8336 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec1/dec4_4/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m1[12] ), .A(\SADR/MAINSADR/oddadd[12] ), .B(
        \SADR/MAINSADR/adrdec1/gcarry[2] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_4/n8327 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec1/dec4_4/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/gg_out[3] ), .A(\SADR/MAINSADR/oddadd[12] ), 
        .B(\SADR/MAINSADR/oddadd[15] ), .C(\SADR/MAINSADR/oddadd[13] ), .D(
        \SADR/MAINSADR/oddadd[14] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec1/dec4_4/U13  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_4/n8331 ), .A(
        \SADR/MAINSADR/adrdec1/dec4_4/n8327 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_4/n8330 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_4/U14  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_4/n8329 ), .A(\SADR/MAINSADR/oddadd[15] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec1/dec4_4/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[15] ), .A(\SADR/MAINSADR/adrdec1/gcarry[2] ), 
        .B(\SADR/MAINSADR/adrdec1/gg_out[3] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_4/n8328 ), .D(
        \SADR/MAINSADR/adrdec1/dec4_4/n8329 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_4/U12  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_4/n8327 ), .A(
        \SADR/MAINSADR/adrdec1/gcarry[2] ), .B(\SADR/MAINSADR/oddadd[12] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec1/dec4_4/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[13] ), .A(
        \SADR/MAINSADR/adrdec1/dec4_4/n8327 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_4/n8330 ), .C(
        \SADR/MAINSADR/adrdec1/dec4_4/n8331 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_4/U15  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_4/n8330 ), .A(\SADR/MAINSADR/oddadd[13] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_4/U11  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_4/n8328 ), .A(\SADR/MAINSADR/oddadd[14] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_4/n8331 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec1/dec4_4/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[14] ), .A(\SADR/MAINSADR/oddadd[14] ), .B(
        \SADR/MAINSADR/adrdec1/dec4_4/n8331 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec1/dec4_6/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m1[20] ), .A(\SADR/MAINSADR/oddadd[20] ), .B(
        \SADR/MAINSADR/adrdec1/gcarry[4] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_6/n8322 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec1/dec4_6/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/dec4_6/gg_out ), .A(\SADR/MAINSADR/oddadd[20] ), 
        .B(\SADR/MAINSADR/oddadd[23] ), .C(\SADR/MAINSADR/oddadd[21] ), .D(
        \SADR/MAINSADR/oddadd[22] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec1/dec4_6/U13  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_6/n8326 ), .A(
        \SADR/MAINSADR/adrdec1/dec4_6/n8322 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_6/n8325 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_6/U14  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_6/n8324 ), .A(\SADR/MAINSADR/oddadd[23] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec1/dec4_6/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[23] ), .A(\SADR/MAINSADR/adrdec1/gcarry[4] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_6/gg_out ), .C(
        \SADR/MAINSADR/adrdec1/dec4_6/n8323 ), .D(
        \SADR/MAINSADR/adrdec1/dec4_6/n8324 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_6/U12  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_6/n8322 ), .A(
        \SADR/MAINSADR/adrdec1/gcarry[4] ), .B(\SADR/MAINSADR/oddadd[20] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec1/dec4_6/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[21] ), .A(
        \SADR/MAINSADR/adrdec1/dec4_6/n8322 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_6/n8325 ), .C(
        \SADR/MAINSADR/adrdec1/dec4_6/n8326 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_6/U15  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_6/n8325 ), .A(\SADR/MAINSADR/oddadd[21] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_6/U11  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_6/n8323 ), .A(\SADR/MAINSADR/oddadd[22] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_6/n8326 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec1/dec4_6/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[22] ), .A(\SADR/MAINSADR/oddadd[22] ), .B(
        \SADR/MAINSADR/adrdec1/dec4_6/n8326 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec1/dec4_5/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m1[16] ), .A(\SADR/MAINSADR/oddadd[16] ), .B(
        \SADR/MAINSADR/adrdec1/gcarry[3] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_5/n8317 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec1/dec4_5/U8  ( .Z(
        \SADR/MAINSADR/adrdec1/gg_out[4] ), .A(\SADR/MAINSADR/oddadd[16] ), 
        .B(\SADR/MAINSADR/oddadd[19] ), .C(\SADR/MAINSADR/oddadd[17] ), .D(
        \SADR/MAINSADR/oddadd[18] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec1/dec4_5/U13  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_5/n8321 ), .A(
        \SADR/MAINSADR/adrdec1/dec4_5/n8317 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_5/n8320 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_5/U14  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_5/n8319 ), .A(\SADR/MAINSADR/oddadd[19] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec1/dec4_5/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[19] ), .A(\SADR/MAINSADR/adrdec1/gcarry[3] ), 
        .B(\SADR/MAINSADR/adrdec1/gg_out[4] ), .C(
        \SADR/MAINSADR/adrdec1/dec4_5/n8318 ), .D(
        \SADR/MAINSADR/adrdec1/dec4_5/n8319 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_5/U12  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_5/n8317 ), .A(
        \SADR/MAINSADR/adrdec1/gcarry[3] ), .B(\SADR/MAINSADR/oddadd[16] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec1/dec4_5/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[17] ), .A(
        \SADR/MAINSADR/adrdec1/dec4_5/n8317 ), .B(
        \SADR/MAINSADR/adrdec1/dec4_5/n8320 ), .C(
        \SADR/MAINSADR/adrdec1/dec4_5/n8321 ) );
    snl_invx05 \SADR/MAINSADR/adrdec1/dec4_5/U15  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_5/n8320 ), .A(\SADR/MAINSADR/oddadd[17] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec1/dec4_5/U11  ( .ZN(
        \SADR/MAINSADR/adrdec1/dec4_5/n8318 ), .A(\SADR/MAINSADR/oddadd[18] ), 
        .B(\SADR/MAINSADR/adrdec1/dec4_5/n8321 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec1/dec4_5/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m1[18] ), .A(\SADR/MAINSADR/oddadd[18] ), .B(
        \SADR/MAINSADR/adrdec1/dec4_5/n8321 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc2/inc4_1/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/gp_out[0] ), .A(\SADR/MAINSADR/oddadd[4] ), .B(
        \SADR/MAINSADR/oddadd[1] ), .C(\SADR/MAINSADR/oddadd[2] ), .D(
        \SADR/MAINSADR/oddadd[3] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_1/U8  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_1/n8314 ), .A(\SADR/MAINSADR/oddadd[1] ), 
        .B(1'b1) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_1/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p2[0] ), .A(\SADR/MAINSADR/oddadd[1] ), .B(1'b1)
         );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_1/U14  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_1/n8316 ), .A(\SADR/MAINSADR/oddadd[3] ), 
        .B(\SADR/MAINSADR/adrinc2/inc4_1/n8315 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc2/inc4_1/U9  ( .Z(
        \SADR/MAINSADR/adrinc2/inc4_1/n8315 ), .A(
        \SADR/MAINSADR/adrinc2/inc4_1/n8314 ), .B(\SADR/MAINSADR/oddadd[2] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_1/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[1] ), .A(\SADR/MAINSADR/oddadd[2] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_1/n8314 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_1/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[3] ), .A(\SADR/MAINSADR/oddadd[4] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_1/n8316 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_1/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p2[2] ), .A(\SADR/MAINSADR/oddadd[3] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_1/n8315 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc2/inc4_2/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/gp_out[1] ), .A(\SADR/MAINSADR/oddadd[8] ), .B(
        \SADR/MAINSADR/oddadd[5] ), .C(\SADR/MAINSADR/oddadd[6] ), .D(
        \SADR/MAINSADR/oddadd[7] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_2/U8  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_2/n8311 ), .A(\SADR/MAINSADR/oddadd[5] ), 
        .B(\SADR/MAINSADR/adrinc2/gp_out[0] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_2/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p2[4] ), .A(\SADR/MAINSADR/oddadd[5] ), .B(
        \SADR/MAINSADR/adrinc2/gp_out[0] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_2/U14  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_2/n8313 ), .A(\SADR/MAINSADR/oddadd[7] ), 
        .B(\SADR/MAINSADR/adrinc2/inc4_2/n8312 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc2/inc4_2/U9  ( .Z(
        \SADR/MAINSADR/adrinc2/inc4_2/n8312 ), .A(
        \SADR/MAINSADR/adrinc2/inc4_2/n8311 ), .B(\SADR/MAINSADR/oddadd[6] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_2/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[5] ), .A(\SADR/MAINSADR/oddadd[6] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_2/n8311 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_2/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[7] ), .A(\SADR/MAINSADR/oddadd[8] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_2/n8313 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_2/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p2[6] ), .A(\SADR/MAINSADR/oddadd[7] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_2/n8312 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc2/inc4_3/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/gp_out[2] ), .A(\SADR/MAINSADR/oddadd[12] ), 
        .B(\SADR/MAINSADR/oddadd[9] ), .C(\SADR/MAINSADR/oddadd[10] ), .D(
        \SADR/MAINSADR/oddadd[11] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_3/U8  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_3/n8308 ), .A(\SADR/MAINSADR/oddadd[9] ), 
        .B(\SADR/MAINSADR/adrinc2/gg_out[1] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_3/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p2[8] ), .A(\SADR/MAINSADR/oddadd[9] ), .B(
        \SADR/MAINSADR/adrinc2/gg_out[1] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_3/U14  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_3/n8310 ), .A(\SADR/MAINSADR/oddadd[11] ), 
        .B(\SADR/MAINSADR/adrinc2/inc4_3/n8309 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc2/inc4_3/U9  ( .Z(
        \SADR/MAINSADR/adrinc2/inc4_3/n8309 ), .A(
        \SADR/MAINSADR/adrinc2/inc4_3/n8308 ), .B(\SADR/MAINSADR/oddadd[10] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_3/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[9] ), .A(\SADR/MAINSADR/oddadd[10] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_3/n8308 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_3/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[11] ), .A(\SADR/MAINSADR/oddadd[12] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_3/n8310 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_3/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p2[10] ), .A(\SADR/MAINSADR/oddadd[11] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_3/n8309 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc2/inc4_4/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/gp_out[3] ), .A(\SADR/MAINSADR/oddadd[16] ), 
        .B(\SADR/MAINSADR/oddadd[13] ), .C(\SADR/MAINSADR/oddadd[14] ), .D(
        \SADR/MAINSADR/oddadd[15] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_4/U8  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_4/n8305 ), .A(\SADR/MAINSADR/oddadd[13] ), 
        .B(\SADR/MAINSADR/adrinc2/gg_out[2] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_4/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p2[12] ), .A(\SADR/MAINSADR/oddadd[13] ), .B(
        \SADR/MAINSADR/adrinc2/gg_out[2] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_4/U14  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_4/n8307 ), .A(\SADR/MAINSADR/oddadd[15] ), 
        .B(\SADR/MAINSADR/adrinc2/inc4_4/n8306 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc2/inc4_4/U9  ( .Z(
        \SADR/MAINSADR/adrinc2/inc4_4/n8306 ), .A(
        \SADR/MAINSADR/adrinc2/inc4_4/n8305 ), .B(\SADR/MAINSADR/oddadd[14] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_4/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[13] ), .A(\SADR/MAINSADR/oddadd[14] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_4/n8305 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_4/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[15] ), .A(\SADR/MAINSADR/oddadd[16] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_4/n8307 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_4/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p2[14] ), .A(\SADR/MAINSADR/oddadd[15] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_4/n8306 ) );
    snl_and04x1 \SADR/MAINSADR/adrinc2/inc4_5/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/gp_out[4] ), .A(\SADR/MAINSADR/oddadd[20] ), 
        .B(\SADR/MAINSADR/oddadd[17] ), .C(\SADR/MAINSADR/oddadd[18] ), .D(
        \SADR/MAINSADR/oddadd[19] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_5/U8  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_5/n8302 ), .A(\SADR/MAINSADR/oddadd[17] ), 
        .B(\SADR/MAINSADR/adrinc2/gg_out[3] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_5/U13  ( .Z(
        \SADR/MAINSADR/oddadd_p2[16] ), .A(\SADR/MAINSADR/oddadd[17] ), .B(
        \SADR/MAINSADR/adrinc2/gg_out[3] ) );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc4_5/U14  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc4_5/n8304 ), .A(\SADR/MAINSADR/oddadd[19] ), 
        .B(\SADR/MAINSADR/adrinc2/inc4_5/n8303 ) );
    snl_and12x1 \SADR/MAINSADR/adrinc2/inc4_5/U9  ( .Z(
        \SADR/MAINSADR/adrinc2/inc4_5/n8303 ), .A(
        \SADR/MAINSADR/adrinc2/inc4_5/n8302 ), .B(\SADR/MAINSADR/oddadd[18] )
         );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_5/U12  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[17] ), .A(\SADR/MAINSADR/oddadd[18] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_5/n8302 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc4_5/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[19] ), .A(\SADR/MAINSADR/oddadd[20] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_5/n8304 ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc4_5/U11  ( .Z(
        \SADR/MAINSADR/oddadd_p2[18] ), .A(\SADR/MAINSADR/oddadd[19] ), .B(
        \SADR/MAINSADR/adrinc2/inc4_5/n8303 ) );
    snl_and03x1 \SADR/MAINSADR/adrinc2/inc3_6/U7  ( .Z(
        \SADR/MAINSADR/adrinc2/inc3_6/gp_out ), .A(\SADR/MAINSADR/oddadd[23] ), 
        .B(\SADR/MAINSADR/oddadd[21] ), .C(\SADR/MAINSADR/oddadd[22] ) );
    snl_and12x1 \SADR/MAINSADR/adrinc2/inc3_6/U8  ( .Z(
        \SADR/MAINSADR/adrinc2/inc3_6/n8300 ), .A(
        \SADR/MAINSADR/adrinc2/inc3_6/n8301 ), .B(\SADR/MAINSADR/oddadd[22] )
         );
    snl_nand02x1 \SADR/MAINSADR/adrinc2/inc3_6/U9  ( .ZN(
        \SADR/MAINSADR/adrinc2/inc3_6/n8301 ), .A(
        \SADR/MAINSADR/adrinc2/gg_out[4] ), .B(\SADR/MAINSADR/oddadd[21] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc3_6/U12  ( .Z(
        \SADR/MAINSADR/oddadd_p2[20] ), .A(\SADR/MAINSADR/adrinc2/gg_out[4] ), 
        .B(\SADR/MAINSADR/oddadd[21] ) );
    snl_xor2x0 \SADR/MAINSADR/adrinc2/inc3_6/U10  ( .Z(
        \SADR/MAINSADR/oddadd_p2[22] ), .A(\SADR/MAINSADR/oddadd[23] ), .B(
        \SADR/MAINSADR/adrinc2/inc3_6/n8300 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrinc2/inc3_6/U11  ( .ZN(
        \SADR/MAINSADR/oddadd_p2[21] ), .A(\SADR/MAINSADR/oddadd[22] ), .B(
        \SADR/MAINSADR/adrinc2/inc3_6/n8301 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec2/dec4_1/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m2[0] ), .A(\SADR/MAINSADR/oddadd[1] ), .B(1'b0), 
        .C(\SADR/MAINSADR/adrdec2/dec4_1/n8294 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec2/dec4_1/U8  ( .Z(
        \SADR/MAINSADR/adrdec2/gg_out[0] ), .A(\SADR/MAINSADR/oddadd[1] ), .B(
        \SADR/MAINSADR/oddadd[4] ), .C(\SADR/MAINSADR/oddadd[2] ), .D(
        \SADR/MAINSADR/oddadd[3] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec2/dec4_1/U13  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_1/n8298 ), .A(
        \SADR/MAINSADR/adrdec2/dec4_1/n8294 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_1/n8297 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_1/U14  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_1/n8296 ), .A(\SADR/MAINSADR/oddadd[4] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec2/dec4_1/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[3] ), .A(1'b0), .B(
        \SADR/MAINSADR/adrdec2/gg_out[0] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_1/n8295 ), .D(
        \SADR/MAINSADR/adrdec2/dec4_1/n8296 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_1/U12  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_1/n8294 ), .A(1'b0), .B(
        \SADR/MAINSADR/oddadd[1] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec2/dec4_1/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[1] ), .A(\SADR/MAINSADR/adrdec2/dec4_1/n8294 
        ), .B(\SADR/MAINSADR/adrdec2/dec4_1/n8297 ), .C(
        \SADR/MAINSADR/adrdec2/dec4_1/n8298 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_1/U15  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_1/n8297 ), .A(\SADR/MAINSADR/oddadd[2] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_1/U11  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_1/n8295 ), .A(\SADR/MAINSADR/oddadd[3] ), 
        .B(\SADR/MAINSADR/adrdec2/dec4_1/n8298 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec2/dec4_1/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[2] ), .A(\SADR/MAINSADR/oddadd[3] ), .B(
        \SADR/MAINSADR/adrdec2/dec4_1/n8298 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec2/dec4_2/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m2[4] ), .A(\SADR/MAINSADR/oddadd[5] ), .B(
        \SADR/MAINSADR/adrdec2/gg_out[0] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_2/n8289 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec2/dec4_2/U8  ( .Z(
        \SADR/MAINSADR/adrdec2/gg_out[1] ), .A(\SADR/MAINSADR/oddadd[5] ), .B(
        \SADR/MAINSADR/oddadd[8] ), .C(\SADR/MAINSADR/oddadd[6] ), .D(
        \SADR/MAINSADR/oddadd[7] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec2/dec4_2/U13  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_2/n8293 ), .A(
        \SADR/MAINSADR/adrdec2/dec4_2/n8289 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_2/n8292 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_2/U14  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_2/n8291 ), .A(\SADR/MAINSADR/oddadd[8] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec2/dec4_2/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[7] ), .A(\SADR/MAINSADR/adrdec2/gg_out[0] ), 
        .B(\SADR/MAINSADR/adrdec2/gg_out[1] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_2/n8290 ), .D(
        \SADR/MAINSADR/adrdec2/dec4_2/n8291 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_2/U12  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_2/n8289 ), .A(
        \SADR/MAINSADR/adrdec2/gg_out[0] ), .B(\SADR/MAINSADR/oddadd[5] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec2/dec4_2/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[5] ), .A(\SADR/MAINSADR/adrdec2/dec4_2/n8289 
        ), .B(\SADR/MAINSADR/adrdec2/dec4_2/n8292 ), .C(
        \SADR/MAINSADR/adrdec2/dec4_2/n8293 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_2/U15  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_2/n8292 ), .A(\SADR/MAINSADR/oddadd[6] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_2/U11  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_2/n8290 ), .A(\SADR/MAINSADR/oddadd[7] ), 
        .B(\SADR/MAINSADR/adrdec2/dec4_2/n8293 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec2/dec4_2/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[6] ), .A(\SADR/MAINSADR/oddadd[7] ), .B(
        \SADR/MAINSADR/adrdec2/dec4_2/n8293 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec2/dec4_3/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m2[8] ), .A(\SADR/MAINSADR/oddadd[9] ), .B(
        \SADR/MAINSADR/adrdec2/gcarry[1] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_3/n8284 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec2/dec4_3/U8  ( .Z(
        \SADR/MAINSADR/adrdec2/gg_out[2] ), .A(\SADR/MAINSADR/oddadd[9] ), .B(
        \SADR/MAINSADR/oddadd[12] ), .C(\SADR/MAINSADR/oddadd[10] ), .D(
        \SADR/MAINSADR/oddadd[11] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec2/dec4_3/U13  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_3/n8288 ), .A(
        \SADR/MAINSADR/adrdec2/dec4_3/n8284 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_3/n8287 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_3/U14  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_3/n8286 ), .A(\SADR/MAINSADR/oddadd[12] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec2/dec4_3/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[11] ), .A(\SADR/MAINSADR/adrdec2/gcarry[1] ), 
        .B(\SADR/MAINSADR/adrdec2/gg_out[2] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_3/n8285 ), .D(
        \SADR/MAINSADR/adrdec2/dec4_3/n8286 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_3/U12  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_3/n8284 ), .A(
        \SADR/MAINSADR/adrdec2/gcarry[1] ), .B(\SADR/MAINSADR/oddadd[9] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec2/dec4_3/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[9] ), .A(\SADR/MAINSADR/adrdec2/dec4_3/n8284 
        ), .B(\SADR/MAINSADR/adrdec2/dec4_3/n8287 ), .C(
        \SADR/MAINSADR/adrdec2/dec4_3/n8288 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_3/U15  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_3/n8287 ), .A(\SADR/MAINSADR/oddadd[10] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_3/U11  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_3/n8285 ), .A(\SADR/MAINSADR/oddadd[11] ), 
        .B(\SADR/MAINSADR/adrdec2/dec4_3/n8288 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec2/dec4_3/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[10] ), .A(\SADR/MAINSADR/oddadd[11] ), .B(
        \SADR/MAINSADR/adrdec2/dec4_3/n8288 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec2/dec4_4/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m2[12] ), .A(\SADR/MAINSADR/oddadd[13] ), .B(
        \SADR/MAINSADR/adrdec2/gcarry[2] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_4/n8279 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec2/dec4_4/U8  ( .Z(
        \SADR/MAINSADR/adrdec2/gg_out[3] ), .A(\SADR/MAINSADR/oddadd[13] ), 
        .B(\SADR/MAINSADR/oddadd[16] ), .C(\SADR/MAINSADR/oddadd[14] ), .D(
        \SADR/MAINSADR/oddadd[15] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec2/dec4_4/U13  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_4/n8283 ), .A(
        \SADR/MAINSADR/adrdec2/dec4_4/n8279 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_4/n8282 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_4/U14  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_4/n8281 ), .A(\SADR/MAINSADR/oddadd[16] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec2/dec4_4/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[15] ), .A(\SADR/MAINSADR/adrdec2/gcarry[2] ), 
        .B(\SADR/MAINSADR/adrdec2/gg_out[3] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_4/n8280 ), .D(
        \SADR/MAINSADR/adrdec2/dec4_4/n8281 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_4/U12  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_4/n8279 ), .A(
        \SADR/MAINSADR/adrdec2/gcarry[2] ), .B(\SADR/MAINSADR/oddadd[13] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec2/dec4_4/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[13] ), .A(
        \SADR/MAINSADR/adrdec2/dec4_4/n8279 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_4/n8282 ), .C(
        \SADR/MAINSADR/adrdec2/dec4_4/n8283 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_4/U15  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_4/n8282 ), .A(\SADR/MAINSADR/oddadd[14] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_4/U11  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_4/n8280 ), .A(\SADR/MAINSADR/oddadd[15] ), 
        .B(\SADR/MAINSADR/adrdec2/dec4_4/n8283 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec2/dec4_4/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[14] ), .A(\SADR/MAINSADR/oddadd[15] ), .B(
        \SADR/MAINSADR/adrdec2/dec4_4/n8283 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec2/dec4_5/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m2[16] ), .A(\SADR/MAINSADR/oddadd[17] ), .B(
        \SADR/MAINSADR/adrdec2/gcarry[3] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_5/n8274 ) );
    snl_or04x1 \SADR/MAINSADR/adrdec2/dec4_5/U8  ( .Z(
        \SADR/MAINSADR/adrdec2/gg_out[4] ), .A(\SADR/MAINSADR/oddadd[17] ), 
        .B(\SADR/MAINSADR/oddadd[20] ), .C(\SADR/MAINSADR/oddadd[18] ), .D(
        \SADR/MAINSADR/oddadd[19] ) );
    snl_nand02x1 \SADR/MAINSADR/adrdec2/dec4_5/U13  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_5/n8278 ), .A(
        \SADR/MAINSADR/adrdec2/dec4_5/n8274 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_5/n8277 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_5/U14  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_5/n8276 ), .A(\SADR/MAINSADR/oddadd[20] )
         );
    snl_oai022x1 \SADR/MAINSADR/adrdec2/dec4_5/U9  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[19] ), .A(\SADR/MAINSADR/adrdec2/gcarry[3] ), 
        .B(\SADR/MAINSADR/adrdec2/gg_out[4] ), .C(
        \SADR/MAINSADR/adrdec2/dec4_5/n8275 ), .D(
        \SADR/MAINSADR/adrdec2/dec4_5/n8276 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_5/U12  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_5/n8274 ), .A(
        \SADR/MAINSADR/adrdec2/gcarry[3] ), .B(\SADR/MAINSADR/oddadd[17] ) );
    snl_oai012x1 \SADR/MAINSADR/adrdec2/dec4_5/U10  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[17] ), .A(
        \SADR/MAINSADR/adrdec2/dec4_5/n8274 ), .B(
        \SADR/MAINSADR/adrdec2/dec4_5/n8277 ), .C(
        \SADR/MAINSADR/adrdec2/dec4_5/n8278 ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec4_5/U15  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_5/n8277 ), .A(\SADR/MAINSADR/oddadd[18] )
         );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec4_5/U11  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec4_5/n8275 ), .A(\SADR/MAINSADR/oddadd[19] ), 
        .B(\SADR/MAINSADR/adrdec2/dec4_5/n8278 ) );
    snl_xnor2x0 \SADR/MAINSADR/adrdec2/dec4_5/U16  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[18] ), .A(\SADR/MAINSADR/oddadd[19] ), .B(
        \SADR/MAINSADR/adrdec2/dec4_5/n8278 ) );
    snl_ao012x1 \SADR/MAINSADR/adrdec2/dec3_6/U7  ( .Z(
        \SADR/MAINSADR/oddadd_m2[20] ), .A(\SADR/MAINSADR/oddadd[21] ), .B(
        \SADR/MAINSADR/adrdec2/gcarry[4] ), .C(
        \SADR/MAINSADR/adrdec2/dec3_6/n8271 ) );
    snl_oai022x1 \SADR/MAINSADR/adrdec2/dec3_6/U8  ( .ZN(
        \SADR/MAINSADR/oddadd_m2[22] ), .A(\SADR/MAINSADR/adrdec2/gcarry[4] ), 
        .B(\SADR/MAINSADR/adrdec2/dec3_6/gg_out ), .C(
        \SADR/MAINSADR/adrdec2/dec3_6/n8272 ), .D(
        \SADR/MAINSADR/adrdec2/dec3_6/n8273 ) );
    snl_xor2x0 \SADR/MAINSADR/adrdec2/dec3_6/U13  ( .Z(
        \SADR/MAINSADR/oddadd_m2[21] ), .A(\SADR/MAINSADR/oddadd[22] ), .B(
        \SADR/MAINSADR/adrdec2/dec3_6/n8271 ) );
    snl_or03x1 \SADR/MAINSADR/adrdec2/dec3_6/U9  ( .Z(
        \SADR/MAINSADR/adrdec2/dec3_6/gg_out ), .A(\SADR/MAINSADR/oddadd[22] ), 
        .B(\SADR/MAINSADR/oddadd[21] ), .C(\SADR/MAINSADR/oddadd[23] ) );
    snl_invx05 \SADR/MAINSADR/adrdec2/dec3_6/U12  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec3_6/n8273 ), .A(\SADR/MAINSADR/oddadd[23] )
         );
    snl_and12x1 \SADR/MAINSADR/adrdec2/dec3_6/U10  ( .Z(
        \SADR/MAINSADR/adrdec2/dec3_6/n8272 ), .A(\SADR/MAINSADR/oddadd[22] ), 
        .B(\SADR/MAINSADR/adrdec2/dec3_6/n8271 ) );
    snl_nor02x1 \SADR/MAINSADR/adrdec2/dec3_6/U11  ( .ZN(
        \SADR/MAINSADR/adrdec2/dec3_6/n8271 ), .A(
        \SADR/MAINSADR/adrdec2/gcarry[4] ), .B(\SADR/MAINSADR/oddadd[21] ) );
    snl_and04x1 \REGF/pbmemff21/pbinc19k_1/inc4_1/U7  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gp_out[0] ), .A(\pk_pc_h[3] ), .B(
        \pk_pc_h[0] ), .C(\pk_pc_h[1] ), .D(\pk_pc_h[2] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_1/U8  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6966 ), .A(\pk_pc_h[0] ), .B(1'b1)
         );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_1/U13  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[0] ), .A(\pk_pc_h[0] ), .B(1'b1) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_1/U14  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6968 ), .A(\pk_pc_h[2] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6967 ) );
    snl_and12x1 \REGF/pbmemff21/pbinc19k_1/inc4_1/U9  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6967 ), .A(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6966 ), .B(\pk_pc_h[1] ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_1/U12  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[1] ), .A(\pk_pc_h[1] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6966 ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_1/U10  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[3] ), .A(\pk_pc_h[3] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6968 ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_1/U11  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[2] ), .A(\pk_pc_h[2] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_1/n6967 ) );
    snl_and03x1 \REGF/pbmemff21/pbinc19k_1/inc3_5/U7  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/inc3_5/gp_out ), .A(\pk_pc_h[18] ), .B(
        \pk_pc_h[16] ), .C(\pk_pc_h[17] ) );
    snl_and12x1 \REGF/pbmemff21/pbinc19k_1/inc3_5/U8  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6964 ), .A(
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6965 ), .B(\pk_pc_h[17] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc3_5/U9  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6965 ), .A(
        \REGF/pbmemff21/pbinc19k_1/gg_out[3] ), .B(\pk_pc_h[16] ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc3_5/U12  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[16] ), .A(
        \REGF/pbmemff21/pbinc19k_1/gg_out[3] ), .B(\pk_pc_h[16] ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc3_5/U10  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[18] ), .A(\pk_pc_h[18] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6964 ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc3_5/U11  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[17] ), .A(\pk_pc_h[17] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc3_5/n6965 ) );
    snl_and04x1 \REGF/pbmemff21/pbinc19k_1/inc4_2/U7  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gp_out[1] ), .A(\pk_pc_h[7] ), .B(
        \pk_pc_h[4] ), .C(\pk_pc_h[5] ), .D(\pk_pc_h[6] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_2/U8  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6961 ), .A(\pk_pc_h[4] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gp_out[0] ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_2/U13  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[4] ), .A(\pk_pc_h[4] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gp_out[0] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_2/U14  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6963 ), .A(\pk_pc_h[6] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6962 ) );
    snl_and12x1 \REGF/pbmemff21/pbinc19k_1/inc4_2/U9  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6962 ), .A(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6961 ), .B(\pk_pc_h[5] ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_2/U12  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[5] ), .A(\pk_pc_h[5] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6961 ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_2/U10  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[7] ), .A(\pk_pc_h[7] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6963 ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_2/U11  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[6] ), .A(\pk_pc_h[6] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_2/n6962 ) );
    snl_and04x1 \REGF/pbmemff21/pbinc19k_1/inc4_3/U7  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gp_out[2] ), .A(\pk_pc_h[11] ), .B(
        \pk_pc_h[8] ), .C(\pk_pc_h[9] ), .D(\pk_pc_h[10] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_3/U8  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6958 ), .A(\pk_pc_h[8] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gg_out[1] ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_3/U13  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[8] ), .A(\pk_pc_h[8] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gg_out[1] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_3/U14  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6960 ), .A(\pk_pc_h[10] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6959 ) );
    snl_and12x1 \REGF/pbmemff21/pbinc19k_1/inc4_3/U9  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6959 ), .A(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6958 ), .B(\pk_pc_h[9] ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_3/U12  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[9] ), .A(\pk_pc_h[9] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6958 ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_3/U10  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[11] ), .A(\pk_pc_h[11] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6960 ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_3/U11  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[10] ), .A(\pk_pc_h[10] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_3/n6959 ) );
    snl_and04x1 \REGF/pbmemff21/pbinc19k_1/inc4_4/U7  ( .Z(
        \REGF/pbmemff21/pbinc19k_1/gp_out[3] ), .A(\pk_pc_h[15] ), .B(
        \pk_pc_h[12] ), .C(\pk_pc_h[13] ), .D(\pk_pc_h[14] ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_4/U8  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6953 ), .A(\pk_pc_h[12] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gg_out[2] ) );
    snl_aoi022x1 \REGF/pbmemff21/pbinc19k_1/inc4_4/U13  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[13] ), .A(\pk_pc_h[13] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6957 ), .C(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6954 ), .D(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6953 ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_4/U14  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[12] ), .A(\pk_pc_h[12] ), .B(
        \REGF/pbmemff21/pbinc19k_1/gg_out[2] ) );
    snl_invx05 \REGF/pbmemff21/pbinc19k_1/inc4_4/U9  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6954 ), .A(\pk_pc_h[13] ) );
    snl_xor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_4/U12  ( .Z(
        \REGF/pbmemff21/RO_PC19BT[14] ), .A(\pk_pc_h[14] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6955 ) );
    snl_nor02x1 \REGF/pbmemff21/pbinc19k_1/inc4_4/U10  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6955 ), .A(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6954 ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6953 ) );
    snl_nand02x1 \REGF/pbmemff21/pbinc19k_1/inc4_4/U15  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6956 ), .A(\pk_pc_h[14] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6955 ) );
    snl_xnor2x0 \REGF/pbmemff21/pbinc19k_1/inc4_4/U11  ( .ZN(
        \REGF/pbmemff21/RO_PC19BT[15] ), .A(\pk_pc_h[15] ), .B(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6956 ) );
    snl_invx05 \REGF/pbmemff21/pbinc19k_1/inc4_4/U16  ( .ZN(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6957 ), .A(
        \REGF/pbmemff21/pbinc19k_1/inc4_4/n6953 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10623 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10624 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10625 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10626 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10623 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10627 ), .D(
        \SADR/ADDIDX/add_w_x/add0/n10628 ), .E(
        \SADR/ADDIDX/add_w_x/add0/n10629 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10639 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10638 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10640 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_x/add0/n10641 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10626 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10642 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10642 ), .A(\pk_indw_h[0] ), .B(
        \pk_indx_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10644 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10623 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10637 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10640 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10626 ), .A(\pk_indw_h[0] ), .B(
        \pk_indx_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10625 ), .A(\pk_indw_h[4] ), .B(
        \pk_indx_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10647 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10648 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10652 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add0/U26  ( .Z(\SADR/pgaddwx[0] ), .A(1'b0
        ), .B(\SADR/ADDIDX/add_w_x/add0/n10641 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_x/gg_out[0] ), .A(\SADR/ADDIDX/add_w_x/add0/n10629 
        ), .B(\SADR/ADDIDX/add_w_x/add0/n10630 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10631 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10635 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10636 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10637 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10638 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10646 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10650 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10626 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10628 ), .D(
        \SADR/ADDIDX/add_w_x/add0/n10651 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10623 ), .A(\pk_indw_h[4] ), .B(
        \pk_indx_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10624 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10646 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10653 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10634 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add0/U20  ( .Z(\SADR/pgaddwx[1] ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10636 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10639 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10648 ), .A(\pk_indw_h[2] ), .B(
        \pk_indx_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10643 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10651 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10627 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10654 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10632 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10631 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10629 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10630 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10643 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10644 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10625 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add0/U17  ( .Z(\SADR/pgaddwx[4] ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10645 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10624 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10628 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10648 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10637 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10640 ), .A(\pk_indw_h[1] ), .B(
        \pk_indx_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10634 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10654 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10638 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10649 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10629 ), .A(\pk_indw_h[5] ), .B(
        \pk_indx_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10636 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10626 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10650 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10642 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10633 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10634 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10627 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add0/U19  ( .Z(\SADR/pgaddwx[2] ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10647 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10635 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_x/add0/n10651 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10642 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10628 ), .C(
        \SADR/ADDIDX/add_w_x/add0/n10648 ), .D(
        \SADR/ADDIDX/add_w_x/add0/n10649 ), .E(
        \SADR/ADDIDX/add_w_x/add0/n10652 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10653 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10627 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add0/U16  ( .Z(\SADR/pgaddwx[5] ), .A(
        \SADR/ADDIDX/add_w_x/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10632 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add0/U18  ( .Z(\SADR/pgaddwx[3] ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10646 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10633 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10627 ), .A(\pk_indw_h[3] ), .B(
        \pk_indx_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_x/add0/n10631 ), .A(\pk_indw_h[5] ), .B(
        \pk_indx_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10649 ), .A(\pk_indw_h[1] ), .B(
        \pk_indx_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10650 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10652 ), .A(\pk_indw_h[2] ), .B(
        \pk_indx_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10654 ), .A(\pk_indw_h[3] ), .B(
        \pk_indx_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x/add0/n10645 ), .A(
        \SADR/ADDIDX/add_w_x/add0/n10644 ), .B(
        \SADR/ADDIDX/add_w_x/add0/n10625 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10591 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10592 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10593 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x/gp_out[1] ), .A(\SADR/ADDIDX/add_w_x/add1/n10594 
        ), .B(\SADR/ADDIDX/add_w_x/add1/n10591 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10595 ), .D(
        \SADR/ADDIDX/add_w_x/add1/n10596 ), .E(
        \SADR/ADDIDX/add_w_x/add1/n10597 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10607 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10606 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10608 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_x/add1/n10609 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10594 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10610 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10610 ), .A(\pk_indw_h[6] ), .B(
        \pk_indx_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10612 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10591 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10605 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10608 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10594 ), .A(\pk_indw_h[6] ), .B(
        \pk_indx_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10593 ), .A(\pk_indw_h[10] ), .B(
        \pk_indx_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10615 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10616 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10620 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add1/U26  ( .Z(\SADR/pgaddwx[6] ), .A(
        \SADR/ADDIDX/add_w_x/gg_out[0] ), .B(\SADR/ADDIDX/add_w_x/add1/n10609 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_x/gg_out[1] ), .A(\SADR/ADDIDX/add_w_x/add1/n10597 
        ), .B(\SADR/ADDIDX/add_w_x/add1/n10598 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10599 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10603 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10604 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10605 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10606 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10614 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10618 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10594 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10596 ), .D(
        \SADR/ADDIDX/add_w_x/add1/n10619 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10591 ), .A(\pk_indw_h[10] ), .B(
        \pk_indx_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10592 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10614 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10621 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10602 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add1/U20  ( .Z(\SADR/pgaddwx[7] ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10604 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10607 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10616 ), .A(\pk_indw_h[8] ), .B(
        \pk_indx_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10611 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10619 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10595 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10622 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10600 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10599 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10597 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10598 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10611 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10612 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10593 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add1/U17  ( .Z(\SADR/pgaddwx[10] ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10613 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10592 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10596 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10616 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10605 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10608 ), .A(\pk_indw_h[7] ), .B(
        \pk_indx_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10602 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10622 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10606 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10617 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10597 ), .A(\pk_indw_h[11] ), .B(
        \pk_indx_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10604 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10594 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10618 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10610 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10601 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10602 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10595 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add1/U19  ( .Z(\SADR/pgaddwx[8] ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10615 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10603 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_x/add1/n10619 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10610 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10596 ), .C(
        \SADR/ADDIDX/add_w_x/add1/n10616 ), .D(
        \SADR/ADDIDX/add_w_x/add1/n10617 ), .E(
        \SADR/ADDIDX/add_w_x/add1/n10620 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10621 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10595 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add1/U16  ( .Z(\SADR/pgaddwx[11] ), .A(
        \SADR/ADDIDX/add_w_x/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10600 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add1/U18  ( .Z(\SADR/pgaddwx[9] ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10614 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10601 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10595 ), .A(\pk_indw_h[9] ), .B(
        \pk_indx_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_x/add1/n10599 ), .A(\pk_indw_h[11] ), .B(
        \pk_indx_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10617 ), .A(\pk_indw_h[7] ), .B(
        \pk_indx_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10618 ), .A(\SADR/ADDIDX/add_w_x/gg_out[0] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10620 ), .A(\pk_indw_h[8] ), .B(
        \pk_indx_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10622 ), .A(\pk_indw_h[9] ), .B(
        \pk_indx_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x/add1/n10613 ), .A(
        \SADR/ADDIDX/add_w_x/add1/n10612 ), .B(
        \SADR/ADDIDX/add_w_x/add1/n10593 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10559 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10560 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10561 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x/gp_out[2] ), .A(\SADR/ADDIDX/add_w_x/add2/n10562 
        ), .B(\SADR/ADDIDX/add_w_x/add2/n10559 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10563 ), .D(
        \SADR/ADDIDX/add_w_x/add2/n10564 ), .E(
        \SADR/ADDIDX/add_w_x/add2/n10565 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10575 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10574 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10576 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_x/add2/n10577 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10562 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10578 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10578 ), .A(\pk_indw_h[12] ), .B(
        \pk_indx_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10580 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10559 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10573 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10576 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10562 ), .A(\pk_indw_h[12] ), .B(
        \pk_indx_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10561 ), .A(\pk_indw_h[16] ), .B(
        \pk_indx_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10583 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10584 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10588 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add2/U26  ( .Z(\SADR/pgaddwx[12] ), .A(
        \SADR/ADDIDX/add_w_x/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10577 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_x/gg_out[2] ), .A(\SADR/ADDIDX/add_w_x/add2/n10565 
        ), .B(\SADR/ADDIDX/add_w_x/add2/n10566 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10567 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10571 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10572 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10573 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10574 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10582 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10586 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10562 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10564 ), .D(
        \SADR/ADDIDX/add_w_x/add2/n10587 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10559 ), .A(\pk_indw_h[16] ), .B(
        \pk_indx_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10560 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10582 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10589 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10570 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add2/U20  ( .Z(\SADR/pgaddwx[13] ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10572 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10575 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10584 ), .A(\pk_indw_h[14] ), .B(
        \pk_indx_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10579 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10587 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10563 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10590 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10568 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10567 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10565 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10566 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10579 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10580 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10561 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add2/U17  ( .Z(\SADR/pgaddwx[16] ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10581 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10560 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10564 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10584 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10573 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10576 ), .A(\pk_indw_h[13] ), .B(
        \pk_indx_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10570 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10590 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10574 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10585 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10565 ), .A(\pk_indw_h[17] ), .B(
        \pk_indx_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10572 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10562 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10586 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10578 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10569 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10570 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10563 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add2/U19  ( .Z(\SADR/pgaddwx[14] ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10583 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10571 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_x/add2/n10587 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10578 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10564 ), .C(
        \SADR/ADDIDX/add_w_x/add2/n10584 ), .D(
        \SADR/ADDIDX/add_w_x/add2/n10585 ), .E(
        \SADR/ADDIDX/add_w_x/add2/n10588 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10589 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10563 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add2/U16  ( .Z(\SADR/pgaddwx[17] ), .A(
        \SADR/ADDIDX/add_w_x/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10568 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add2/U18  ( .Z(\SADR/pgaddwx[15] ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10582 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10569 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10563 ), .A(\pk_indw_h[15] ), .B(
        \pk_indx_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_x/add2/n10567 ), .A(\pk_indw_h[17] ), .B(
        \pk_indx_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10585 ), .A(\pk_indw_h[13] ), .B(
        \pk_indx_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10586 ), .A(
        \SADR/ADDIDX/add_w_x/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10588 ), .A(\pk_indw_h[14] ), .B(
        \pk_indx_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10590 ), .A(\pk_indw_h[15] ), .B(
        \pk_indx_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x/add2/n10581 ), .A(
        \SADR/ADDIDX/add_w_x/add2/n10580 ), .B(
        \SADR/ADDIDX/add_w_x/add2/n10561 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x/c_last ), .A(\SADR/ADDIDX/add_w_x/add3/n10527 ), 
        .B(\SADR/ADDIDX/add_w_x/add3/n10528 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10529 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x/gp_out[3] ), .A(\SADR/ADDIDX/add_w_x/add3/n10530 
        ), .B(\SADR/ADDIDX/add_w_x/add3/n10527 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10531 ), .D(
        \SADR/ADDIDX/add_w_x/add3/n10532 ), .E(
        \SADR/ADDIDX/add_w_x/add3/n10533 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10543 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10542 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10544 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_x/add3/n10545 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10530 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10546 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10546 ), .A(\pk_indw_h[18] ), .B(
        \pk_indx_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10548 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10527 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10541 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10544 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10530 ), .A(\pk_indw_h[18] ), .B(
        \pk_indx_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10529 ), .A(\pk_indw_h[22] ), .B(
        \pk_indx_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10551 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10552 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10556 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add3/U26  ( .Z(\SADR/pgaddwx[18] ), .A(
        \SADR/ADDIDX/add_w_x/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10545 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_x/gg_out[3] ), .A(\SADR/ADDIDX/add_w_x/add3/n10533 
        ), .B(\SADR/ADDIDX/add_w_x/add3/n10534 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10535 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10539 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10540 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10541 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10542 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10550 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10554 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10530 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10532 ), .D(
        \SADR/ADDIDX/add_w_x/add3/n10555 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10527 ), .A(\pk_indw_h[22] ), .B(
        \pk_indx_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10528 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10550 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10557 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10538 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add3/U20  ( .Z(\SADR/pgaddwx[19] ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10540 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10543 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10552 ), .A(\pk_indw_h[20] ), .B(
        \pk_indx_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10547 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10555 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10531 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10558 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10536 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10535 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10533 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10534 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10547 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10548 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10529 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add3/U17  ( .Z(\SADR/pgaddwx[22] ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10549 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10528 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10532 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10552 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10541 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10544 ), .A(\pk_indw_h[19] ), .B(
        \pk_indx_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10538 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10558 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10542 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10553 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10533 ), .A(\pk_indw_h[23] ), .B(
        \pk_indx_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10540 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10530 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10554 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10546 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10537 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10538 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10531 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add3/U19  ( .Z(\SADR/pgaddwx[20] ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10551 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10539 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_x/add3/n10555 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10546 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10532 ), .C(
        \SADR/ADDIDX/add_w_x/add3/n10552 ), .D(
        \SADR/ADDIDX/add_w_x/add3/n10553 ), .E(
        \SADR/ADDIDX/add_w_x/add3/n10556 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10557 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10531 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add3/U16  ( .Z(\SADR/pgaddwx[23] ), .A(
        \SADR/ADDIDX/add_w_x/c_last ), .B(\SADR/ADDIDX/add_w_x/add3/n10536 )
         );
    snl_xor2x0 \SADR/ADDIDX/add_w_x/add3/U18  ( .Z(\SADR/pgaddwx[21] ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10550 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10537 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10531 ), .A(\pk_indw_h[21] ), .B(
        \pk_indx_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_x/add3/n10535 ), .A(\pk_indw_h[23] ), .B(
        \pk_indx_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10553 ), .A(\pk_indw_h[19] ), .B(
        \pk_indx_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10554 ), .A(
        \SADR/ADDIDX/add_w_x/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10556 ), .A(\pk_indw_h[20] ), .B(
        \pk_indx_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10558 ), .A(\pk_indw_h[21] ), .B(
        \pk_indx_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x/add3/n10549 ), .A(
        \SADR/ADDIDX/add_w_x/add3/n10548 ), .B(
        \SADR/ADDIDX/add_w_x/add3/n10529 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10494 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10495 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10496 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10497 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10494 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10498 ), .D(
        \SADR/ADDIDX/add_x_z/add0/n10499 ), .E(
        \SADR/ADDIDX/add_x_z/add0/n10500 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10510 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10509 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10511 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_x_z/add0/n10512 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10497 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10513 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10513 ), .A(\pk_indx_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10515 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10494 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10508 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10511 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10497 ), .A(\pk_indx_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10496 ), .A(\pk_indx_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10518 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10519 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10523 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add0/U26  ( .Z(\SADR/pgaddxz[0] ), .A(1'b0
        ), .B(\SADR/ADDIDX/add_x_z/add0/n10512 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_x_z/gg_out[0] ), .A(\SADR/ADDIDX/add_x_z/add0/n10500 
        ), .B(\SADR/ADDIDX/add_x_z/add0/n10501 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10502 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10506 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10507 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10508 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10509 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10517 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10521 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10497 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10499 ), .D(
        \SADR/ADDIDX/add_x_z/add0/n10522 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10494 ), .A(\pk_indx_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10495 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10517 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10524 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10505 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add0/U20  ( .Z(\SADR/pgaddxz[1] ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10507 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10510 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10519 ), .A(\pk_indx_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10514 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10522 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10498 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10525 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10503 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10502 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10500 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10501 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10514 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10515 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10496 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add0/U17  ( .Z(\SADR/pgaddxz[4] ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10516 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10495 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10499 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10519 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10508 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10511 ), .A(\pk_indx_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10505 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10525 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10509 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10520 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10500 ), .A(\pk_indx_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10507 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10497 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10521 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10513 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10504 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10505 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10498 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add0/U19  ( .Z(\SADR/pgaddxz[2] ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10518 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10506 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_x_z/add0/n10522 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10513 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10499 ), .C(
        \SADR/ADDIDX/add_x_z/add0/n10519 ), .D(
        \SADR/ADDIDX/add_x_z/add0/n10520 ), .E(
        \SADR/ADDIDX/add_x_z/add0/n10523 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10524 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10498 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add0/U16  ( .Z(\SADR/pgaddxz[5] ), .A(
        \SADR/ADDIDX/add_x_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10503 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add0/U18  ( .Z(\SADR/pgaddxz[3] ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10517 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10504 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10498 ), .A(\pk_indx_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_x_z/add0/n10502 ), .A(\pk_indx_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10520 ), .A(\pk_indx_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10521 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10523 ), .A(\pk_indx_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10525 ), .A(\pk_indx_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_x_z/add0/n10516 ), .A(
        \SADR/ADDIDX/add_x_z/add0/n10515 ), .B(
        \SADR/ADDIDX/add_x_z/add0/n10496 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10462 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10463 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10464 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_x_z/gp_out[1] ), .A(\SADR/ADDIDX/add_x_z/add1/n10465 
        ), .B(\SADR/ADDIDX/add_x_z/add1/n10462 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10466 ), .D(
        \SADR/ADDIDX/add_x_z/add1/n10467 ), .E(
        \SADR/ADDIDX/add_x_z/add1/n10468 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10478 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10477 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10479 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_x_z/add1/n10480 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10465 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10481 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10481 ), .A(\pk_indx_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10483 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10462 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10476 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10479 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10465 ), .A(\pk_indx_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10464 ), .A(\pk_indx_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10486 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10487 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10491 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add1/U26  ( .Z(\SADR/pgaddxz[6] ), .A(
        \SADR/ADDIDX/add_x_z/gg_out[0] ), .B(\SADR/ADDIDX/add_x_z/add1/n10480 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_x_z/gg_out[1] ), .A(\SADR/ADDIDX/add_x_z/add1/n10468 
        ), .B(\SADR/ADDIDX/add_x_z/add1/n10469 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10470 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10474 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10475 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10476 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10477 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10485 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10489 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10465 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10467 ), .D(
        \SADR/ADDIDX/add_x_z/add1/n10490 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10462 ), .A(\pk_indx_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10463 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10485 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10492 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10473 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add1/U20  ( .Z(\SADR/pgaddxz[7] ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10475 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10478 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10487 ), .A(\pk_indx_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10482 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10490 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10466 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10493 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10471 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10470 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10468 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10469 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10482 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10483 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10464 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add1/U17  ( .Z(\SADR/pgaddxz[10] ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10484 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10463 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10467 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10487 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10476 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10479 ), .A(\pk_indx_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10473 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10493 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10477 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10488 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10468 ), .A(\pk_indx_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10475 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10465 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10489 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10481 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10472 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10473 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10466 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add1/U19  ( .Z(\SADR/pgaddxz[8] ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10486 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10474 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_x_z/add1/n10490 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10481 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10467 ), .C(
        \SADR/ADDIDX/add_x_z/add1/n10487 ), .D(
        \SADR/ADDIDX/add_x_z/add1/n10488 ), .E(
        \SADR/ADDIDX/add_x_z/add1/n10491 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10492 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10466 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add1/U16  ( .Z(\SADR/pgaddxz[11] ), .A(
        \SADR/ADDIDX/add_x_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10471 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add1/U18  ( .Z(\SADR/pgaddxz[9] ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10485 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10472 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10466 ), .A(\pk_indx_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_x_z/add1/n10470 ), .A(\pk_indx_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10488 ), .A(\pk_indx_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10489 ), .A(\SADR/ADDIDX/add_x_z/gg_out[0] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10491 ), .A(\pk_indx_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10493 ), .A(\pk_indx_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_x_z/add1/n10484 ), .A(
        \SADR/ADDIDX/add_x_z/add1/n10483 ), .B(
        \SADR/ADDIDX/add_x_z/add1/n10464 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10430 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10431 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10432 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_x_z/gp_out[2] ), .A(\SADR/ADDIDX/add_x_z/add2/n10433 
        ), .B(\SADR/ADDIDX/add_x_z/add2/n10430 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10434 ), .D(
        \SADR/ADDIDX/add_x_z/add2/n10435 ), .E(
        \SADR/ADDIDX/add_x_z/add2/n10436 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10446 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10445 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10447 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_x_z/add2/n10448 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10433 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10449 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10449 ), .A(\pk_indx_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10451 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10430 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10444 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10447 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10433 ), .A(\pk_indx_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10432 ), .A(\pk_indx_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10454 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10455 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10459 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add2/U26  ( .Z(\SADR/pgaddxz[12] ), .A(
        \SADR/ADDIDX/add_x_z/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10448 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_x_z/gg_out[2] ), .A(\SADR/ADDIDX/add_x_z/add2/n10436 
        ), .B(\SADR/ADDIDX/add_x_z/add2/n10437 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10438 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10442 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10443 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10444 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10445 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10453 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10457 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10433 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10435 ), .D(
        \SADR/ADDIDX/add_x_z/add2/n10458 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10430 ), .A(\pk_indx_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10431 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10453 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10460 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10441 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add2/U20  ( .Z(\SADR/pgaddxz[13] ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10443 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10446 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10455 ), .A(\pk_indx_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10450 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10458 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10434 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10461 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10439 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10438 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10436 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10437 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10450 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10451 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10432 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add2/U17  ( .Z(\SADR/pgaddxz[16] ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10452 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10431 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10435 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10455 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10444 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10447 ), .A(\pk_indx_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10441 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10461 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10445 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10456 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10436 ), .A(\pk_indx_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10443 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10433 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10457 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10449 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10440 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10441 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10434 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add2/U19  ( .Z(\SADR/pgaddxz[14] ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10454 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10442 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_x_z/add2/n10458 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10449 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10435 ), .C(
        \SADR/ADDIDX/add_x_z/add2/n10455 ), .D(
        \SADR/ADDIDX/add_x_z/add2/n10456 ), .E(
        \SADR/ADDIDX/add_x_z/add2/n10459 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10460 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10434 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add2/U16  ( .Z(\SADR/pgaddxz[17] ), .A(
        \SADR/ADDIDX/add_x_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10439 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add2/U18  ( .Z(\SADR/pgaddxz[15] ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10453 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10440 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10434 ), .A(\pk_indx_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_x_z/add2/n10438 ), .A(\pk_indx_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10456 ), .A(\pk_indx_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10457 ), .A(
        \SADR/ADDIDX/add_x_z/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10459 ), .A(\pk_indx_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10461 ), .A(\pk_indx_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_x_z/add2/n10452 ), .A(
        \SADR/ADDIDX/add_x_z/add2/n10451 ), .B(
        \SADR/ADDIDX/add_x_z/add2/n10432 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_x_z/c_last ), .A(\SADR/ADDIDX/add_x_z/add3/n10398 ), 
        .B(\SADR/ADDIDX/add_x_z/add3/n10399 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10400 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_x_z/gp_out[3] ), .A(\SADR/ADDIDX/add_x_z/add3/n10401 
        ), .B(\SADR/ADDIDX/add_x_z/add3/n10398 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10402 ), .D(
        \SADR/ADDIDX/add_x_z/add3/n10403 ), .E(
        \SADR/ADDIDX/add_x_z/add3/n10404 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10414 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10413 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10415 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_x_z/add3/n10416 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10401 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10417 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10417 ), .A(\pk_indx_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10419 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10398 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10412 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10415 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10401 ), .A(\pk_indx_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10400 ), .A(\pk_indx_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10422 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10423 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10427 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add3/U26  ( .Z(\SADR/pgaddxz[18] ), .A(
        \SADR/ADDIDX/add_x_z/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10416 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_x_z/gg_out[3] ), .A(\SADR/ADDIDX/add_x_z/add3/n10404 
        ), .B(\SADR/ADDIDX/add_x_z/add3/n10405 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10406 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10410 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10411 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10412 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10413 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10421 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10425 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10401 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10403 ), .D(
        \SADR/ADDIDX/add_x_z/add3/n10426 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10398 ), .A(\pk_indx_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10399 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10421 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10428 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10409 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add3/U20  ( .Z(\SADR/pgaddxz[19] ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10411 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10414 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10423 ), .A(\pk_indx_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10418 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10426 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10402 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10429 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10407 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10406 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10404 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10405 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10418 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10419 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10400 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add3/U17  ( .Z(\SADR/pgaddxz[22] ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10420 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10399 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10403 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10423 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10412 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10415 ), .A(\pk_indx_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10409 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10429 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10413 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10424 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10404 ), .A(\pk_indx_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10411 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10401 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10425 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10417 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10408 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10409 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10402 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add3/U19  ( .Z(\SADR/pgaddxz[20] ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10422 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10410 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_x_z/add3/n10426 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10417 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10403 ), .C(
        \SADR/ADDIDX/add_x_z/add3/n10423 ), .D(
        \SADR/ADDIDX/add_x_z/add3/n10424 ), .E(
        \SADR/ADDIDX/add_x_z/add3/n10427 ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10428 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10402 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add3/U16  ( .Z(\SADR/pgaddxz[23] ), .A(
        \SADR/ADDIDX/add_x_z/c_last ), .B(\SADR/ADDIDX/add_x_z/add3/n10407 )
         );
    snl_xor2x0 \SADR/ADDIDX/add_x_z/add3/U18  ( .Z(\SADR/pgaddxz[21] ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10421 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10408 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10402 ), .A(\pk_indx_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_x_z/add3/n10406 ), .A(\pk_indx_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10424 ), .A(\pk_indx_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_x_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10425 ), .A(
        \SADR/ADDIDX/add_x_z/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10427 ), .A(\pk_indx_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10429 ), .A(\pk_indx_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_x_z/add3/n10420 ), .A(
        \SADR/ADDIDX/add_x_z/add3/n10419 ), .B(
        \SADR/ADDIDX/add_x_z/add3/n10400 ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10365 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10366 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10367 ) );
    snl_nor05x1 \SADR/ADDIDX/add_y_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10368 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10365 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10369 ), .D(
        \SADR/ADDIDX/add_y_z/add0/n10370 ), .E(
        \SADR/ADDIDX/add_y_z/add0/n10371 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10381 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10380 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10382 ) );
    snl_and12x1 \SADR/ADDIDX/add_y_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_y_z/add0/n10383 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10368 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10384 ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10384 ), .A(\pk_indy_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10386 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10365 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10379 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10382 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10368 ), .A(\pk_indy_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10367 ), .A(\pk_indy_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10389 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10390 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10394 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add0/U26  ( .Z(\SADR/pgaddyz[0] ), .A(1'b0
        ), .B(\SADR/ADDIDX/add_y_z/add0/n10383 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_y_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_y_z/gg_out[0] ), .A(\SADR/ADDIDX/add_y_z/add0/n10371 
        ), .B(\SADR/ADDIDX/add_y_z/add0/n10372 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10373 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10377 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10378 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10379 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10380 ) );
    snl_oai013x0 \SADR/ADDIDX/add_y_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10388 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10392 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10368 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10370 ), .D(
        \SADR/ADDIDX/add_y_z/add0/n10393 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10365 ), .A(\pk_indy_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10366 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10388 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10395 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10376 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add0/U20  ( .Z(\SADR/pgaddyz[1] ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10378 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10381 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10390 ), .A(\pk_indy_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10385 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10393 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10369 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10396 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10374 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10373 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10371 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_y_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10372 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10385 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10386 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10367 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add0/U17  ( .Z(\SADR/pgaddyz[4] ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10387 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10366 ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10370 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10390 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10379 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10382 ), .A(\pk_indy_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10376 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10396 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10380 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10391 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10371 ), .A(\pk_indy_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10378 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10368 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10392 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10384 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10375 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10376 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10369 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add0/U19  ( .Z(\SADR/pgaddyz[2] ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10389 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10377 ) );
    snl_oa122x1 \SADR/ADDIDX/add_y_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_y_z/add0/n10393 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10384 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10370 ), .C(
        \SADR/ADDIDX/add_y_z/add0/n10390 ), .D(
        \SADR/ADDIDX/add_y_z/add0/n10391 ), .E(
        \SADR/ADDIDX/add_y_z/add0/n10394 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10395 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10369 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add0/U16  ( .Z(\SADR/pgaddyz[5] ), .A(
        \SADR/ADDIDX/add_y_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10374 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add0/U18  ( .Z(\SADR/pgaddyz[3] ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10388 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10375 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10369 ), .A(\pk_indy_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_y_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_y_z/add0/n10373 ), .A(\pk_indy_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10391 ), .A(\pk_indy_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10392 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10394 ), .A(\pk_indy_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10396 ), .A(\pk_indy_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_y_z/add0/n10387 ), .A(
        \SADR/ADDIDX/add_y_z/add0/n10386 ), .B(
        \SADR/ADDIDX/add_y_z/add0/n10367 ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10333 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10334 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10335 ) );
    snl_nor05x1 \SADR/ADDIDX/add_y_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_y_z/gp_out[1] ), .A(\SADR/ADDIDX/add_y_z/add1/n10336 
        ), .B(\SADR/ADDIDX/add_y_z/add1/n10333 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10337 ), .D(
        \SADR/ADDIDX/add_y_z/add1/n10338 ), .E(
        \SADR/ADDIDX/add_y_z/add1/n10339 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10349 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10348 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10350 ) );
    snl_and12x1 \SADR/ADDIDX/add_y_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_y_z/add1/n10351 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10336 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10352 ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10352 ), .A(\pk_indy_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10354 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10333 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10347 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10350 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10336 ), .A(\pk_indy_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10335 ), .A(\pk_indy_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10357 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10358 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10362 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add1/U26  ( .Z(\SADR/pgaddyz[6] ), .A(
        \SADR/ADDIDX/add_y_z/gg_out[0] ), .B(\SADR/ADDIDX/add_y_z/add1/n10351 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_y_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_y_z/gg_out[1] ), .A(\SADR/ADDIDX/add_y_z/add1/n10339 
        ), .B(\SADR/ADDIDX/add_y_z/add1/n10340 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10341 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10345 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10346 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10347 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10348 ) );
    snl_oai013x0 \SADR/ADDIDX/add_y_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10356 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10360 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10336 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10338 ), .D(
        \SADR/ADDIDX/add_y_z/add1/n10361 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10333 ), .A(\pk_indy_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10334 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10356 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10363 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10344 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add1/U20  ( .Z(\SADR/pgaddyz[7] ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10346 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10349 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10358 ), .A(\pk_indy_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10353 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10361 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10337 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10364 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10342 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10341 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10339 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_y_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10340 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10353 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10354 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10335 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add1/U17  ( .Z(\SADR/pgaddyz[10] ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10355 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10334 ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10338 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10358 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10347 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10350 ), .A(\pk_indy_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10344 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10364 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10348 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10359 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10339 ), .A(\pk_indy_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10346 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10336 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10360 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10352 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10343 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10344 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10337 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add1/U19  ( .Z(\SADR/pgaddyz[8] ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10357 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10345 ) );
    snl_oa122x1 \SADR/ADDIDX/add_y_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_y_z/add1/n10361 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10352 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10338 ), .C(
        \SADR/ADDIDX/add_y_z/add1/n10358 ), .D(
        \SADR/ADDIDX/add_y_z/add1/n10359 ), .E(
        \SADR/ADDIDX/add_y_z/add1/n10362 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10363 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10337 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add1/U16  ( .Z(\SADR/pgaddyz[11] ), .A(
        \SADR/ADDIDX/add_y_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10342 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add1/U18  ( .Z(\SADR/pgaddyz[9] ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10356 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10343 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10337 ), .A(\pk_indy_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_y_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_y_z/add1/n10341 ), .A(\pk_indy_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10359 ), .A(\pk_indy_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10360 ), .A(\SADR/ADDIDX/add_y_z/gg_out[0] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10362 ), .A(\pk_indy_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10364 ), .A(\pk_indy_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_y_z/add1/n10355 ), .A(
        \SADR/ADDIDX/add_y_z/add1/n10354 ), .B(
        \SADR/ADDIDX/add_y_z/add1/n10335 ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10301 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10302 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10303 ) );
    snl_nor05x1 \SADR/ADDIDX/add_y_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_y_z/gp_out[2] ), .A(\SADR/ADDIDX/add_y_z/add2/n10304 
        ), .B(\SADR/ADDIDX/add_y_z/add2/n10301 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10305 ), .D(
        \SADR/ADDIDX/add_y_z/add2/n10306 ), .E(
        \SADR/ADDIDX/add_y_z/add2/n10307 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10317 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10316 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10318 ) );
    snl_and12x1 \SADR/ADDIDX/add_y_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_y_z/add2/n10319 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10304 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10320 ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10320 ), .A(\pk_indy_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10322 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10301 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10315 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10318 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10304 ), .A(\pk_indy_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10303 ), .A(\pk_indy_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10325 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10326 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10330 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add2/U26  ( .Z(\SADR/pgaddyz[12] ), .A(
        \SADR/ADDIDX/add_y_z/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10319 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_y_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_y_z/gg_out[2] ), .A(\SADR/ADDIDX/add_y_z/add2/n10307 
        ), .B(\SADR/ADDIDX/add_y_z/add2/n10308 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10309 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10313 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10314 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10315 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10316 ) );
    snl_oai013x0 \SADR/ADDIDX/add_y_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10324 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10328 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10304 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10306 ), .D(
        \SADR/ADDIDX/add_y_z/add2/n10329 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10301 ), .A(\pk_indy_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10302 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10324 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10331 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10312 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add2/U20  ( .Z(\SADR/pgaddyz[13] ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10314 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10317 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10326 ), .A(\pk_indy_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10321 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10329 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10305 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10332 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10310 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10309 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10307 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_y_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10308 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10321 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10322 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10303 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add2/U17  ( .Z(\SADR/pgaddyz[16] ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10323 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10302 ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10306 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10326 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10315 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10318 ), .A(\pk_indy_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10312 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10332 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10316 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10327 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10307 ), .A(\pk_indy_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10314 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10304 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10328 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10320 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10311 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10312 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10305 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add2/U19  ( .Z(\SADR/pgaddyz[14] ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10325 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10313 ) );
    snl_oa122x1 \SADR/ADDIDX/add_y_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_y_z/add2/n10329 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10320 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10306 ), .C(
        \SADR/ADDIDX/add_y_z/add2/n10326 ), .D(
        \SADR/ADDIDX/add_y_z/add2/n10327 ), .E(
        \SADR/ADDIDX/add_y_z/add2/n10330 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10331 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10305 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add2/U16  ( .Z(\SADR/pgaddyz[17] ), .A(
        \SADR/ADDIDX/add_y_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10310 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add2/U18  ( .Z(\SADR/pgaddyz[15] ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10324 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10311 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10305 ), .A(\pk_indy_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_y_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_y_z/add2/n10309 ), .A(\pk_indy_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10327 ), .A(\pk_indy_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10328 ), .A(
        \SADR/ADDIDX/add_y_z/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10330 ), .A(\pk_indy_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10332 ), .A(\pk_indy_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_y_z/add2/n10323 ), .A(
        \SADR/ADDIDX/add_y_z/add2/n10322 ), .B(
        \SADR/ADDIDX/add_y_z/add2/n10303 ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_y_z/c_last ), .A(\SADR/ADDIDX/add_y_z/add3/n10269 ), 
        .B(\SADR/ADDIDX/add_y_z/add3/n10270 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10271 ) );
    snl_nor05x1 \SADR/ADDIDX/add_y_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_y_z/gp_out[3] ), .A(\SADR/ADDIDX/add_y_z/add3/n10272 
        ), .B(\SADR/ADDIDX/add_y_z/add3/n10269 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10273 ), .D(
        \SADR/ADDIDX/add_y_z/add3/n10274 ), .E(
        \SADR/ADDIDX/add_y_z/add3/n10275 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10285 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10284 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10286 ) );
    snl_and12x1 \SADR/ADDIDX/add_y_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_y_z/add3/n10287 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10272 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10288 ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10288 ), .A(\pk_indy_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10290 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10269 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10283 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10286 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10272 ), .A(\pk_indy_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10271 ), .A(\pk_indy_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10293 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10294 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10298 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add3/U26  ( .Z(\SADR/pgaddyz[18] ), .A(
        \SADR/ADDIDX/add_y_z/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10287 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_y_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_y_z/gg_out[3] ), .A(\SADR/ADDIDX/add_y_z/add3/n10275 
        ), .B(\SADR/ADDIDX/add_y_z/add3/n10276 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10277 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10281 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10282 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10283 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10284 ) );
    snl_oai013x0 \SADR/ADDIDX/add_y_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10292 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10296 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10272 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10274 ), .D(
        \SADR/ADDIDX/add_y_z/add3/n10297 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10269 ), .A(\pk_indy_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_y_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10270 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10292 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10299 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10280 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add3/U20  ( .Z(\SADR/pgaddyz[19] ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10282 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10285 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10294 ), .A(\pk_indy_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10289 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10297 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10273 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10300 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10278 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10277 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10275 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_y_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10276 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10289 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10290 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10271 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add3/U17  ( .Z(\SADR/pgaddyz[22] ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10291 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10270 ) );
    snl_nand12x1 \SADR/ADDIDX/add_y_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10274 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10294 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10283 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10286 ), .A(\pk_indy_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10280 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10300 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10284 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10295 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10275 ), .A(\pk_indy_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_y_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10282 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10272 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10296 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10288 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10279 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10280 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10273 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add3/U19  ( .Z(\SADR/pgaddyz[20] ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10293 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10281 ) );
    snl_oa122x1 \SADR/ADDIDX/add_y_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_y_z/add3/n10297 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10288 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10274 ), .C(
        \SADR/ADDIDX/add_y_z/add3/n10294 ), .D(
        \SADR/ADDIDX/add_y_z/add3/n10295 ), .E(
        \SADR/ADDIDX/add_y_z/add3/n10298 ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10299 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10273 ) );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add3/U16  ( .Z(\SADR/pgaddyz[23] ), .A(
        \SADR/ADDIDX/add_y_z/c_last ), .B(\SADR/ADDIDX/add_y_z/add3/n10278 )
         );
    snl_xor2x0 \SADR/ADDIDX/add_y_z/add3/U18  ( .Z(\SADR/pgaddyz[21] ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10292 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10279 ) );
    snl_nor02x1 \SADR/ADDIDX/add_y_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10273 ), .A(\pk_indy_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_y_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_y_z/add3/n10277 ), .A(\pk_indy_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10295 ), .A(\pk_indy_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_y_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10296 ), .A(
        \SADR/ADDIDX/add_y_z/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10298 ), .A(\pk_indy_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10300 ), .A(\pk_indy_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_y_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_y_z/add3/n10291 ), .A(
        \SADR/ADDIDX/add_y_z/add3/n10290 ), .B(
        \SADR/ADDIDX/add_y_z/add3/n10271 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10236 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10237 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10238 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10239 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10236 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10240 ), .D(
        \SADR/ADDIDX/add_w_y/add0/n10241 ), .E(
        \SADR/ADDIDX/add_w_y/add0/n10242 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10252 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10251 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10253 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_y/add0/n10254 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10239 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10255 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10255 ), .A(\pk_indw_h[0] ), .B(
        \pk_indy_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10257 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10236 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10250 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10253 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10239 ), .A(\pk_indw_h[0] ), .B(
        \pk_indy_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10238 ), .A(\pk_indw_h[4] ), .B(
        \pk_indy_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10260 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10261 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10265 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add0/U26  ( .Z(\SADR/pgaddwy[0] ), .A(1'b0
        ), .B(\SADR/ADDIDX/add_w_y/add0/n10254 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_y/gg_out[0] ), .A(\SADR/ADDIDX/add_w_y/add0/n10242 
        ), .B(\SADR/ADDIDX/add_w_y/add0/n10243 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10244 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10248 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10249 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10250 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10251 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10259 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10263 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10239 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10241 ), .D(
        \SADR/ADDIDX/add_w_y/add0/n10264 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10236 ), .A(\pk_indw_h[4] ), .B(
        \pk_indy_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10237 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10259 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10266 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10247 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add0/U20  ( .Z(\SADR/pgaddwy[1] ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10249 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10252 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10261 ), .A(\pk_indw_h[2] ), .B(
        \pk_indy_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10256 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10264 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10240 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10267 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10245 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10244 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10242 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10243 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10256 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10257 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10238 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add0/U17  ( .Z(\SADR/pgaddwy[4] ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10258 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10237 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10241 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10261 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10250 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10253 ), .A(\pk_indw_h[1] ), .B(
        \pk_indy_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10247 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10267 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10251 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10262 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10242 ), .A(\pk_indw_h[5] ), .B(
        \pk_indy_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10249 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10239 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10263 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10255 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10246 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10247 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10240 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add0/U19  ( .Z(\SADR/pgaddwy[2] ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10260 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10248 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_y/add0/n10264 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10255 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10241 ), .C(
        \SADR/ADDIDX/add_w_y/add0/n10261 ), .D(
        \SADR/ADDIDX/add_w_y/add0/n10262 ), .E(
        \SADR/ADDIDX/add_w_y/add0/n10265 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10266 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10240 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add0/U16  ( .Z(\SADR/pgaddwy[5] ), .A(
        \SADR/ADDIDX/add_w_y/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10245 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add0/U18  ( .Z(\SADR/pgaddwy[3] ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10259 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10246 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10240 ), .A(\pk_indw_h[3] ), .B(
        \pk_indy_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_y/add0/n10244 ), .A(\pk_indw_h[5] ), .B(
        \pk_indy_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10262 ), .A(\pk_indw_h[1] ), .B(
        \pk_indy_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10263 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10265 ), .A(\pk_indw_h[2] ), .B(
        \pk_indy_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10267 ), .A(\pk_indw_h[3] ), .B(
        \pk_indy_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y/add0/n10258 ), .A(
        \SADR/ADDIDX/add_w_y/add0/n10257 ), .B(
        \SADR/ADDIDX/add_w_y/add0/n10238 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10204 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10205 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10206 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y/gp_out[1] ), .A(\SADR/ADDIDX/add_w_y/add1/n10207 
        ), .B(\SADR/ADDIDX/add_w_y/add1/n10204 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10208 ), .D(
        \SADR/ADDIDX/add_w_y/add1/n10209 ), .E(
        \SADR/ADDIDX/add_w_y/add1/n10210 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10220 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10219 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10221 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_y/add1/n10222 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10207 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10223 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10223 ), .A(\pk_indw_h[6] ), .B(
        \pk_indy_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10225 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10204 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10218 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10221 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10207 ), .A(\pk_indw_h[6] ), .B(
        \pk_indy_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10206 ), .A(\pk_indw_h[10] ), .B(
        \pk_indy_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10228 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10229 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10233 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add1/U26  ( .Z(\SADR/pgaddwy[6] ), .A(
        \SADR/ADDIDX/add_w_y/gg_out[0] ), .B(\SADR/ADDIDX/add_w_y/add1/n10222 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_y/gg_out[1] ), .A(\SADR/ADDIDX/add_w_y/add1/n10210 
        ), .B(\SADR/ADDIDX/add_w_y/add1/n10211 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10212 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10216 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10217 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10218 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10219 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10227 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10231 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10207 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10209 ), .D(
        \SADR/ADDIDX/add_w_y/add1/n10232 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10204 ), .A(\pk_indw_h[10] ), .B(
        \pk_indy_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10205 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10227 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10234 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10215 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add1/U20  ( .Z(\SADR/pgaddwy[7] ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10217 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10220 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10229 ), .A(\pk_indw_h[8] ), .B(
        \pk_indy_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10224 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10232 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10208 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10235 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10213 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10212 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10210 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10211 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10224 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10225 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10206 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add1/U17  ( .Z(\SADR/pgaddwy[10] ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10226 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10205 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10209 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10229 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10218 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10221 ), .A(\pk_indw_h[7] ), .B(
        \pk_indy_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10215 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10235 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10219 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10230 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10210 ), .A(\pk_indw_h[11] ), .B(
        \pk_indy_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10217 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10207 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10231 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10223 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10214 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10215 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10208 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add1/U19  ( .Z(\SADR/pgaddwy[8] ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10228 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10216 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_y/add1/n10232 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10223 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10209 ), .C(
        \SADR/ADDIDX/add_w_y/add1/n10229 ), .D(
        \SADR/ADDIDX/add_w_y/add1/n10230 ), .E(
        \SADR/ADDIDX/add_w_y/add1/n10233 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10234 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10208 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add1/U16  ( .Z(\SADR/pgaddwy[11] ), .A(
        \SADR/ADDIDX/add_w_y/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10213 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add1/U18  ( .Z(\SADR/pgaddwy[9] ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10227 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10214 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10208 ), .A(\pk_indw_h[9] ), .B(
        \pk_indy_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_y/add1/n10212 ), .A(\pk_indw_h[11] ), .B(
        \pk_indy_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10230 ), .A(\pk_indw_h[7] ), .B(
        \pk_indy_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10231 ), .A(\SADR/ADDIDX/add_w_y/gg_out[0] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10233 ), .A(\pk_indw_h[8] ), .B(
        \pk_indy_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10235 ), .A(\pk_indw_h[9] ), .B(
        \pk_indy_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y/add1/n10226 ), .A(
        \SADR/ADDIDX/add_w_y/add1/n10225 ), .B(
        \SADR/ADDIDX/add_w_y/add1/n10206 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10172 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10173 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10174 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y/gp_out[2] ), .A(\SADR/ADDIDX/add_w_y/add2/n10175 
        ), .B(\SADR/ADDIDX/add_w_y/add2/n10172 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10176 ), .D(
        \SADR/ADDIDX/add_w_y/add2/n10177 ), .E(
        \SADR/ADDIDX/add_w_y/add2/n10178 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10188 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10187 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10189 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_y/add2/n10190 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10175 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10191 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10191 ), .A(\pk_indw_h[12] ), .B(
        \pk_indy_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10193 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10172 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10186 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10189 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10175 ), .A(\pk_indw_h[12] ), .B(
        \pk_indy_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10174 ), .A(\pk_indw_h[16] ), .B(
        \pk_indy_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10196 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10197 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10201 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add2/U26  ( .Z(\SADR/pgaddwy[12] ), .A(
        \SADR/ADDIDX/add_w_y/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10190 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_y/gg_out[2] ), .A(\SADR/ADDIDX/add_w_y/add2/n10178 
        ), .B(\SADR/ADDIDX/add_w_y/add2/n10179 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10180 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10184 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10185 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10186 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10187 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10195 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10199 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10175 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10177 ), .D(
        \SADR/ADDIDX/add_w_y/add2/n10200 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10172 ), .A(\pk_indw_h[16] ), .B(
        \pk_indy_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10173 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10195 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10202 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10183 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add2/U20  ( .Z(\SADR/pgaddwy[13] ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10185 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10188 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10197 ), .A(\pk_indw_h[14] ), .B(
        \pk_indy_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10192 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10200 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10176 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10203 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10181 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10180 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10178 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10179 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10192 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10193 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10174 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add2/U17  ( .Z(\SADR/pgaddwy[16] ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10194 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10173 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10177 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10197 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10186 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10189 ), .A(\pk_indw_h[13] ), .B(
        \pk_indy_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10183 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10203 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10187 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10198 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10178 ), .A(\pk_indw_h[17] ), .B(
        \pk_indy_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10185 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10175 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10199 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10191 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10182 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10183 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10176 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add2/U19  ( .Z(\SADR/pgaddwy[14] ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10196 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10184 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_y/add2/n10200 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10191 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10177 ), .C(
        \SADR/ADDIDX/add_w_y/add2/n10197 ), .D(
        \SADR/ADDIDX/add_w_y/add2/n10198 ), .E(
        \SADR/ADDIDX/add_w_y/add2/n10201 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10202 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10176 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add2/U16  ( .Z(\SADR/pgaddwy[17] ), .A(
        \SADR/ADDIDX/add_w_y/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10181 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add2/U18  ( .Z(\SADR/pgaddwy[15] ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10195 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10182 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10176 ), .A(\pk_indw_h[15] ), .B(
        \pk_indy_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_y/add2/n10180 ), .A(\pk_indw_h[17] ), .B(
        \pk_indy_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10198 ), .A(\pk_indw_h[13] ), .B(
        \pk_indy_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10199 ), .A(
        \SADR/ADDIDX/add_w_y/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10201 ), .A(\pk_indw_h[14] ), .B(
        \pk_indy_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10203 ), .A(\pk_indw_h[15] ), .B(
        \pk_indy_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y/add2/n10194 ), .A(
        \SADR/ADDIDX/add_w_y/add2/n10193 ), .B(
        \SADR/ADDIDX/add_w_y/add2/n10174 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y/c_last ), .A(\SADR/ADDIDX/add_w_y/add3/n10140 ), 
        .B(\SADR/ADDIDX/add_w_y/add3/n10141 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10142 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y/gp_out[3] ), .A(\SADR/ADDIDX/add_w_y/add3/n10143 
        ), .B(\SADR/ADDIDX/add_w_y/add3/n10140 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10144 ), .D(
        \SADR/ADDIDX/add_w_y/add3/n10145 ), .E(
        \SADR/ADDIDX/add_w_y/add3/n10146 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10156 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10155 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10157 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_y/add3/n10158 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10143 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10159 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10159 ), .A(\pk_indw_h[18] ), .B(
        \pk_indy_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10161 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10140 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10154 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10157 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10143 ), .A(\pk_indw_h[18] ), .B(
        \pk_indy_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10142 ), .A(\pk_indw_h[22] ), .B(
        \pk_indy_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10164 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10165 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10169 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add3/U26  ( .Z(\SADR/pgaddwy[18] ), .A(
        \SADR/ADDIDX/add_w_y/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10158 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_y/gg_out[3] ), .A(\SADR/ADDIDX/add_w_y/add3/n10146 
        ), .B(\SADR/ADDIDX/add_w_y/add3/n10147 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10148 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10152 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10153 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10154 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10155 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10163 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10167 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10143 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10145 ), .D(
        \SADR/ADDIDX/add_w_y/add3/n10168 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10140 ), .A(\pk_indw_h[22] ), .B(
        \pk_indy_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10141 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10163 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10170 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10151 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add3/U20  ( .Z(\SADR/pgaddwy[19] ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10153 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10156 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10165 ), .A(\pk_indw_h[20] ), .B(
        \pk_indy_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10160 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10168 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10144 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10171 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10149 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10148 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10146 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10147 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10160 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10161 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10142 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add3/U17  ( .Z(\SADR/pgaddwy[22] ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10162 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10141 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10145 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10165 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10154 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10157 ), .A(\pk_indw_h[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10151 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10171 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10155 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10166 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10146 ), .A(\pk_indw_h[23] ), .B(
        \pk_indy_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10153 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10143 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10167 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10159 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10150 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10151 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10144 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add3/U19  ( .Z(\SADR/pgaddwy[20] ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10164 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10152 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_y/add3/n10168 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10159 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10145 ), .C(
        \SADR/ADDIDX/add_w_y/add3/n10165 ), .D(
        \SADR/ADDIDX/add_w_y/add3/n10166 ), .E(
        \SADR/ADDIDX/add_w_y/add3/n10169 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10170 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10144 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add3/U16  ( .Z(\SADR/pgaddwy[23] ), .A(
        \SADR/ADDIDX/add_w_y/c_last ), .B(\SADR/ADDIDX/add_w_y/add3/n10149 )
         );
    snl_xor2x0 \SADR/ADDIDX/add_w_y/add3/U18  ( .Z(\SADR/pgaddwy[21] ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10163 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10150 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10144 ), .A(\pk_indw_h[21] ), .B(
        \pk_indy_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_y/add3/n10148 ), .A(\pk_indw_h[23] ), .B(
        \pk_indy_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10166 ), .A(\pk_indw_h[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10167 ), .A(
        \SADR/ADDIDX/add_w_y/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10169 ), .A(\pk_indw_h[20] ), .B(
        \pk_indy_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10171 ), .A(\pk_indw_h[21] ), .B(
        \pk_indy_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y/add3/n10162 ), .A(
        \SADR/ADDIDX/add_w_y/add3/n10161 ), .B(
        \SADR/ADDIDX/add_w_y/add3/n10142 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10107 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10108 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10109 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10110 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10107 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10111 ), .D(
        \SADR/ADDIDX/add_w_x_y/add0/n10112 ), .E(
        \SADR/ADDIDX/add_w_x_y/add0/n10113 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10123 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10122 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10124 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add0/n10125 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10110 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10126 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10126 ), .A(\SADR/pgaddwx[0] ), .B(
        \pk_indy_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10128 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10107 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10121 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10124 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10110 ), .A(\SADR/pgaddwx[0] ), .B(
        \pk_indy_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10109 ), .A(\SADR/pgaddwx[4] ), .B(
        \pk_indy_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10131 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10132 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10136 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add0/U26  ( .Z(\SADR/pgaddwxy[0] ), .A(
        1'b0), .B(\SADR/ADDIDX/add_w_x_y/add0/n10125 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y/gg_out[0] ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10113 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10114 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10115 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10119 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10120 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10121 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10122 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10130 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10134 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10110 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10112 ), .D(
        \SADR/ADDIDX/add_w_x_y/add0/n10135 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10107 ), .A(\SADR/pgaddwx[4] ), .B(
        \pk_indy_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10108 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10130 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10137 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10118 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add0/U20  ( .Z(\SADR/pgaddwxy[1] ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10120 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10123 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10132 ), .A(\SADR/pgaddwx[2] ), .B(
        \pk_indy_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10127 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10135 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10111 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10138 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10116 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10115 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10113 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10114 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10127 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10128 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10109 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add0/U17  ( .Z(\SADR/pgaddwxy[4] ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10129 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10108 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10112 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10132 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10121 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10124 ), .A(\SADR/pgaddwx[1] ), .B(
        \pk_indy_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10118 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10138 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10122 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10133 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10113 ), .A(\SADR/pgaddwx[5] ), .B(
        \pk_indy_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10120 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10110 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10134 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10126 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10117 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10118 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10111 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add0/U19  ( .Z(\SADR/pgaddwxy[2] ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10131 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10119 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add0/n10135 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10126 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10112 ), .C(
        \SADR/ADDIDX/add_w_x_y/add0/n10132 ), .D(
        \SADR/ADDIDX/add_w_x_y/add0/n10133 ), .E(
        \SADR/ADDIDX/add_w_x_y/add0/n10136 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10137 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10111 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add0/U16  ( .Z(\SADR/pgaddwxy[5] ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10116 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add0/U18  ( .Z(\SADR/pgaddwxy[3] ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10130 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10117 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10111 ), .A(\SADR/pgaddwx[3] ), .B(
        \pk_indy_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add0/n10115 ), .A(\SADR/pgaddwx[5] ), .B(
        \pk_indy_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10133 ), .A(\SADR/pgaddwx[1] ), .B(
        \pk_indy_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10134 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10136 ), .A(\SADR/pgaddwx[2] ), .B(
        \pk_indy_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10138 ), .A(\SADR/pgaddwx[3] ), .B(
        \pk_indy_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add0/n10129 ), .A(
        \SADR/ADDIDX/add_w_x_y/add0/n10128 ), .B(
        \SADR/ADDIDX/add_w_x_y/add0/n10109 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10075 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10076 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10077 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/gp_out[1] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10078 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10075 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10079 ), .D(
        \SADR/ADDIDX/add_w_x_y/add1/n10080 ), .E(
        \SADR/ADDIDX/add_w_x_y/add1/n10081 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10091 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10090 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10092 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add1/n10093 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10078 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10094 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10094 ), .A(\SADR/pgaddwx[6] ), .B(
        \pk_indy_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10096 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10075 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10089 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10092 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10078 ), .A(\SADR/pgaddwx[6] ), .B(
        \pk_indy_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10077 ), .A(\SADR/pgaddwx[10] ), .B(
        \pk_indy_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10099 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10100 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10104 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add1/U26  ( .Z(\SADR/pgaddwxy[6] ), .A(
        \SADR/ADDIDX/add_w_x_y/gg_out[0] ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10093 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y/gg_out[1] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10081 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10082 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10083 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10087 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10088 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10089 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10090 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10098 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10102 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10078 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10080 ), .D(
        \SADR/ADDIDX/add_w_x_y/add1/n10103 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10075 ), .A(\SADR/pgaddwx[10] ), .B(
        \pk_indy_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10076 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10098 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10105 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10086 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add1/U20  ( .Z(\SADR/pgaddwxy[7] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10088 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10091 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10100 ), .A(\SADR/pgaddwx[8] ), .B(
        \pk_indy_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10095 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10103 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10079 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10106 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10084 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10083 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10081 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10082 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10095 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10096 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10077 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add1/U17  ( .Z(\SADR/pgaddwxy[10] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10097 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10076 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10080 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10100 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10089 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10092 ), .A(\SADR/pgaddwx[7] ), .B(
        \pk_indy_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10086 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10106 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10090 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10101 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10081 ), .A(\SADR/pgaddwx[11] ), .B(
        \pk_indy_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10088 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10078 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10102 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10094 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10085 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10086 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10079 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add1/U19  ( .Z(\SADR/pgaddwxy[8] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10099 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10087 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add1/n10103 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10094 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10080 ), .C(
        \SADR/ADDIDX/add_w_x_y/add1/n10100 ), .D(
        \SADR/ADDIDX/add_w_x_y/add1/n10101 ), .E(
        \SADR/ADDIDX/add_w_x_y/add1/n10104 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10105 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10079 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add1/U16  ( .Z(\SADR/pgaddwxy[11] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10084 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add1/U18  ( .Z(\SADR/pgaddwxy[9] ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10098 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10085 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10079 ), .A(\SADR/pgaddwx[9] ), .B(
        \pk_indy_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add1/n10083 ), .A(\SADR/pgaddwx[11] ), .B(
        \pk_indy_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10101 ), .A(\SADR/pgaddwx[7] ), .B(
        \pk_indy_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10102 ), .A(
        \SADR/ADDIDX/add_w_x_y/gg_out[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10104 ), .A(\SADR/pgaddwx[8] ), .B(
        \pk_indy_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10106 ), .A(\SADR/pgaddwx[9] ), .B(
        \pk_indy_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add1/n10097 ), .A(
        \SADR/ADDIDX/add_w_x_y/add1/n10096 ), .B(
        \SADR/ADDIDX/add_w_x_y/add1/n10077 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10043 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10044 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10045 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/gp_out[2] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10046 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10043 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10047 ), .D(
        \SADR/ADDIDX/add_w_x_y/add2/n10048 ), .E(
        \SADR/ADDIDX/add_w_x_y/add2/n10049 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10059 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10058 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10060 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add2/n10061 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10046 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10062 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10062 ), .A(\SADR/pgaddwx[12] ), .B(
        \pk_indy_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10064 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10043 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10057 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10060 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10046 ), .A(\SADR/pgaddwx[12] ), .B(
        \pk_indy_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10045 ), .A(\SADR/pgaddwx[16] ), .B(
        \pk_indy_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10067 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10068 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10072 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add2/U26  ( .Z(\SADR/pgaddwxy[12] ), .A(
        \SADR/ADDIDX/add_w_x_y/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10061 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y/gg_out[2] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10049 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10050 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10051 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10055 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10056 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10057 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10058 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10066 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10070 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10046 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10048 ), .D(
        \SADR/ADDIDX/add_w_x_y/add2/n10071 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10043 ), .A(\SADR/pgaddwx[16] ), .B(
        \pk_indy_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10044 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10066 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10073 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10054 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add2/U20  ( .Z(\SADR/pgaddwxy[13] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10056 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10059 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10068 ), .A(\SADR/pgaddwx[14] ), .B(
        \pk_indy_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10063 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10071 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10047 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10074 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10052 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10051 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10049 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10050 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10063 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10064 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10045 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add2/U17  ( .Z(\SADR/pgaddwxy[16] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10065 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10044 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10048 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10068 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10057 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10060 ), .A(\SADR/pgaddwx[13] ), .B(
        \pk_indy_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10054 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10074 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10058 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10069 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10049 ), .A(\SADR/pgaddwx[17] ), .B(
        \pk_indy_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10056 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10046 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10070 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10062 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10053 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10054 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10047 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add2/U19  ( .Z(\SADR/pgaddwxy[14] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10067 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10055 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add2/n10071 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10062 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10048 ), .C(
        \SADR/ADDIDX/add_w_x_y/add2/n10068 ), .D(
        \SADR/ADDIDX/add_w_x_y/add2/n10069 ), .E(
        \SADR/ADDIDX/add_w_x_y/add2/n10072 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10073 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10047 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add2/U16  ( .Z(\SADR/pgaddwxy[17] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10052 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add2/U18  ( .Z(\SADR/pgaddwxy[15] ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10066 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10053 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10047 ), .A(\SADR/pgaddwx[15] ), .B(
        \pk_indy_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add2/n10051 ), .A(\SADR/pgaddwx[17] ), .B(
        \pk_indy_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10069 ), .A(\SADR/pgaddwx[13] ), .B(
        \pk_indy_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10070 ), .A(
        \SADR/ADDIDX/add_w_x_y/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10072 ), .A(\SADR/pgaddwx[14] ), .B(
        \pk_indy_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10074 ), .A(\SADR/pgaddwx[15] ), .B(
        \pk_indy_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add2/n10065 ), .A(
        \SADR/ADDIDX/add_w_x_y/add2/n10064 ), .B(
        \SADR/ADDIDX/add_w_x_y/add2/n10045 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10011 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10012 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10013 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/gp_out[3] ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10014 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10011 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10015 ), .D(
        \SADR/ADDIDX/add_w_x_y/add3/n10016 ), .E(
        \SADR/ADDIDX/add_w_x_y/add3/n10017 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10027 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10026 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10028 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add3/n10029 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10014 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10030 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10030 ), .A(\SADR/pgaddwx[18] ), .B(
        \pk_indy_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10032 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10011 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10025 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10028 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10014 ), .A(\SADR/pgaddwx[18] ), .B(
        \pk_indy_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10013 ), .A(\SADR/pgaddwx[22] ), .B(
        \pk_indy_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10035 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10036 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10040 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add3/U26  ( .Z(\SADR/pgaddwxy[18] ), .A(
        \SADR/ADDIDX/add_w_x_y/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10029 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y/gg_out[3] ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10017 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10018 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10019 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10023 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10024 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10025 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10026 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10034 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10038 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10014 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10016 ), .D(
        \SADR/ADDIDX/add_w_x_y/add3/n10039 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10011 ), .A(\SADR/pgaddwx[22] ), .B(
        \pk_indy_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10012 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10034 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10041 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10022 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add3/U20  ( .Z(\SADR/pgaddwxy[19] ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10024 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10027 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10036 ), .A(\SADR/pgaddwx[20] ), .B(
        \pk_indy_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10031 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10039 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10015 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10042 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10020 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10019 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10017 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10018 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10031 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10032 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10013 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add3/U17  ( .Z(\SADR/pgaddwxy[22] ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10033 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10012 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10016 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10036 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10025 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10028 ), .A(\SADR/pgaddwx[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10022 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10042 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10026 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10037 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10017 ), .A(\SADR/pgaddwx[23] ), .B(
        \pk_indy_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10024 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10014 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10038 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10030 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10021 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10022 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10015 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add3/U19  ( .Z(\SADR/pgaddwxy[20] ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10035 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10023 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add3/n10039 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10030 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10016 ), .C(
        \SADR/ADDIDX/add_w_x_y/add3/n10036 ), .D(
        \SADR/ADDIDX/add_w_x_y/add3/n10037 ), .E(
        \SADR/ADDIDX/add_w_x_y/add3/n10040 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10041 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10015 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add3/U16  ( .Z(\SADR/pgaddwxy[23] ), .A(
        \SADR/ADDIDX/add_w_x_y/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10020 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y/add3/U18  ( .Z(\SADR/pgaddwxy[21] ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10034 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10021 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10015 ), .A(\SADR/pgaddwx[21] ), .B(
        \pk_indy_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y/add3/n10019 ), .A(\SADR/pgaddwx[23] ), .B(
        \pk_indy_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10037 ), .A(\SADR/pgaddwx[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10038 ), .A(
        \SADR/ADDIDX/add_w_x_y/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10040 ), .A(\SADR/pgaddwx[20] ), .B(
        \pk_indy_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10042 ), .A(\SADR/pgaddwx[21] ), .B(
        \pk_indy_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y/add3/n10033 ), .A(
        \SADR/ADDIDX/add_w_x_y/add3/n10032 ), .B(
        \SADR/ADDIDX/add_w_x_y/add3/n10013 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9978 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9979 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9980 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9981 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9978 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9982 ), .D(
        \SADR/ADDIDX/add_x_y_z/add0/n9983 ), .E(
        \SADR/ADDIDX/add_x_y_z/add0/n9984 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9994 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9993 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9995 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add0/n9996 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9981 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9997 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9997 ), .A(\SADR/pgaddyz[0] ), .B(
        \pk_indx_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9999 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9978 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9992 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9995 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9981 ), .A(\SADR/pgaddyz[0] ), .B(
        \pk_indx_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9980 ), .A(\SADR/pgaddyz[4] ), .B(
        \pk_indx_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10002 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10003 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n10007 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add0/U26  ( .Z(\SADR/pgaddxyz[0] ), .A(
        1'b0), .B(\SADR/ADDIDX/add_x_y_z/add0/n9996 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_x_y_z/gg_out[0] ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9984 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9985 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9986 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9990 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9991 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9992 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9993 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10001 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10005 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9981 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9983 ), .D(
        \SADR/ADDIDX/add_x_y_z/add0/n10006 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9978 ), .A(\SADR/pgaddyz[4] ), .B(
        \pk_indx_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9979 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10001 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n10008 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9989 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add0/U20  ( .Z(\SADR/pgaddxyz[1] ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9991 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9994 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10003 ), .A(\SADR/pgaddyz[2] ), .B(
        \pk_indx_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9998 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10006 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9982 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n10009 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9987 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9986 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9984 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9985 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9998 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9999 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9980 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add0/U17  ( .Z(\SADR/pgaddxyz[4] ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10000 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9979 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9983 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10003 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9992 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9995 ), .A(\SADR/pgaddyz[1] ), .B(
        \pk_indx_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9989 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10009 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9993 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10004 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9984 ), .A(\SADR/pgaddyz[5] ), .B(
        \pk_indx_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9991 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9981 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n10005 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n9997 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9988 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9989 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9982 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add0/U19  ( .Z(\SADR/pgaddxyz[2] ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10002 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9990 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add0/n10006 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9997 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9983 ), .C(
        \SADR/ADDIDX/add_x_y_z/add0/n10003 ), .D(
        \SADR/ADDIDX/add_x_y_z/add0/n10004 ), .E(
        \SADR/ADDIDX/add_x_y_z/add0/n10007 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10008 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9982 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add0/U16  ( .Z(\SADR/pgaddxyz[5] ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9987 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add0/U18  ( .Z(\SADR/pgaddxyz[3] ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n10001 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9988 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n9982 ), .A(\SADR/pgaddyz[3] ), .B(
        \pk_indx_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add0/n9986 ), .A(\SADR/pgaddyz[5] ), .B(
        \pk_indx_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10004 ), .A(\SADR/pgaddyz[1] ), .B(
        \pk_indx_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10005 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10007 ), .A(\SADR/pgaddyz[2] ), .B(
        \pk_indx_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10009 ), .A(\SADR/pgaddyz[3] ), .B(
        \pk_indx_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add0/n10000 ), .A(
        \SADR/ADDIDX/add_x_y_z/add0/n9999 ), .B(
        \SADR/ADDIDX/add_x_y_z/add0/n9980 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9946 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9947 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9948 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/gp_out[1] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9949 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9946 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9950 ), .D(
        \SADR/ADDIDX/add_x_y_z/add1/n9951 ), .E(
        \SADR/ADDIDX/add_x_y_z/add1/n9952 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9962 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9961 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9963 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add1/n9964 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9949 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9965 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9965 ), .A(\SADR/pgaddyz[6] ), .B(
        \pk_indx_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9967 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9946 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9960 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9963 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9949 ), .A(\SADR/pgaddyz[6] ), .B(
        \pk_indx_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9948 ), .A(\SADR/pgaddyz[10] ), .B(
        \pk_indx_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9970 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9971 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9975 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add1/U26  ( .Z(\SADR/pgaddxyz[6] ), .A(
        \SADR/ADDIDX/add_x_y_z/gg_out[0] ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9964 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_x_y_z/gg_out[1] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9952 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9953 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9954 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9958 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9959 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9960 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9961 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9969 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9973 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9949 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9951 ), .D(
        \SADR/ADDIDX/add_x_y_z/add1/n9974 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9946 ), .A(\SADR/pgaddyz[10] ), .B(
        \pk_indx_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9947 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9969 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9976 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9957 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add1/U20  ( .Z(\SADR/pgaddxyz[7] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9959 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9962 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9971 ), .A(\SADR/pgaddyz[8] ), .B(
        \pk_indx_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9966 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9974 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9950 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9977 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9955 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9954 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9952 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9953 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9966 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9967 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9948 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add1/U17  ( .Z(\SADR/pgaddxyz[10] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9968 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9947 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9951 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9971 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9960 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9963 ), .A(\SADR/pgaddyz[7] ), .B(
        \pk_indx_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9957 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9977 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9961 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9972 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9952 ), .A(\SADR/pgaddyz[11] ), .B(
        \pk_indx_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9959 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9949 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9973 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9965 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9956 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9957 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9950 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add1/U19  ( .Z(\SADR/pgaddxyz[8] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9970 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9958 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add1/n9974 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9965 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9951 ), .C(
        \SADR/ADDIDX/add_x_y_z/add1/n9971 ), .D(
        \SADR/ADDIDX/add_x_y_z/add1/n9972 ), .E(
        \SADR/ADDIDX/add_x_y_z/add1/n9975 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9976 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9950 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add1/U16  ( .Z(\SADR/pgaddxyz[11] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9955 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add1/U18  ( .Z(\SADR/pgaddxyz[9] ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9969 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9956 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9950 ), .A(\SADR/pgaddyz[9] ), .B(
        \pk_indx_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add1/n9954 ), .A(\SADR/pgaddyz[11] ), .B(
        \pk_indx_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9972 ), .A(\SADR/pgaddyz[7] ), .B(
        \pk_indx_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9973 ), .A(
        \SADR/ADDIDX/add_x_y_z/gg_out[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9975 ), .A(\SADR/pgaddyz[8] ), .B(
        \pk_indx_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9977 ), .A(\SADR/pgaddyz[9] ), .B(
        \pk_indx_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add1/n9968 ), .A(
        \SADR/ADDIDX/add_x_y_z/add1/n9967 ), .B(
        \SADR/ADDIDX/add_x_y_z/add1/n9948 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9914 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9915 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9916 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/gp_out[2] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9917 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9914 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9918 ), .D(
        \SADR/ADDIDX/add_x_y_z/add2/n9919 ), .E(
        \SADR/ADDIDX/add_x_y_z/add2/n9920 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9930 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9929 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9931 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add2/n9932 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9917 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9933 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9933 ), .A(\SADR/pgaddyz[12] ), .B(
        \pk_indx_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9935 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9914 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9928 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9931 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9917 ), .A(\SADR/pgaddyz[12] ), .B(
        \pk_indx_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9916 ), .A(\SADR/pgaddyz[16] ), .B(
        \pk_indx_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9938 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9939 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9943 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add2/U26  ( .Z(\SADR/pgaddxyz[12] ), .A(
        \SADR/ADDIDX/add_x_y_z/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9932 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_x_y_z/gg_out[2] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9920 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9921 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9922 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9926 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9927 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9928 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9929 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9937 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9941 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9917 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9919 ), .D(
        \SADR/ADDIDX/add_x_y_z/add2/n9942 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9914 ), .A(\SADR/pgaddyz[16] ), .B(
        \pk_indx_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9915 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9937 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9944 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9925 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add2/U20  ( .Z(\SADR/pgaddxyz[13] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9927 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9930 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9939 ), .A(\SADR/pgaddyz[14] ), .B(
        \pk_indx_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9934 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9942 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9918 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9945 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9923 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9922 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9920 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9921 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9934 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9935 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9916 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add2/U17  ( .Z(\SADR/pgaddxyz[16] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9936 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9915 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9919 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9939 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9928 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9931 ), .A(\SADR/pgaddyz[13] ), .B(
        \pk_indx_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9925 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9945 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9929 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9940 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9920 ), .A(\SADR/pgaddyz[17] ), .B(
        \pk_indx_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9927 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9917 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9941 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9933 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9924 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9925 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9918 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add2/U19  ( .Z(\SADR/pgaddxyz[14] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9938 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9926 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add2/n9942 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9933 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9919 ), .C(
        \SADR/ADDIDX/add_x_y_z/add2/n9939 ), .D(
        \SADR/ADDIDX/add_x_y_z/add2/n9940 ), .E(
        \SADR/ADDIDX/add_x_y_z/add2/n9943 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9944 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9918 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add2/U16  ( .Z(\SADR/pgaddxyz[17] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9923 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add2/U18  ( .Z(\SADR/pgaddxyz[15] ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9937 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9924 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9918 ), .A(\SADR/pgaddyz[15] ), .B(
        \pk_indx_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add2/n9922 ), .A(\SADR/pgaddyz[17] ), .B(
        \pk_indx_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9940 ), .A(\SADR/pgaddyz[13] ), .B(
        \pk_indx_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9941 ), .A(
        \SADR/ADDIDX/add_x_y_z/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9943 ), .A(\SADR/pgaddyz[14] ), .B(
        \pk_indx_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9945 ), .A(\SADR/pgaddyz[15] ), .B(
        \pk_indx_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add2/n9936 ), .A(
        \SADR/ADDIDX/add_x_y_z/add2/n9935 ), .B(
        \SADR/ADDIDX/add_x_y_z/add2/n9916 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/c_last ), .A(\SADR/ADDIDX/add_x_y_z/add3/n9882 
        ), .B(\SADR/ADDIDX/add_x_y_z/add3/n9883 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9884 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/gp_out[3] ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9885 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9882 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9886 ), .D(
        \SADR/ADDIDX/add_x_y_z/add3/n9887 ), .E(
        \SADR/ADDIDX/add_x_y_z/add3/n9888 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9898 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9897 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9899 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add3/n9900 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9885 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9901 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9901 ), .A(\SADR/pgaddyz[18] ), .B(
        \pk_indx_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9903 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9882 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9896 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9899 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9885 ), .A(\SADR/pgaddyz[18] ), .B(
        \pk_indx_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9884 ), .A(\SADR/pgaddyz[22] ), .B(
        \pk_indx_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9906 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9907 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9911 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add3/U26  ( .Z(\SADR/pgaddxyz[18] ), .A(
        \SADR/ADDIDX/add_x_y_z/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9900 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_x_y_z/gg_out[3] ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9888 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9889 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9890 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9894 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9895 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9896 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9897 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9905 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9909 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9885 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9887 ), .D(
        \SADR/ADDIDX/add_x_y_z/add3/n9910 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9882 ), .A(\SADR/pgaddyz[22] ), .B(
        \pk_indx_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9883 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9905 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9912 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9893 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add3/U20  ( .Z(\SADR/pgaddxyz[19] ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9895 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9898 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9907 ), .A(\SADR/pgaddyz[20] ), .B(
        \pk_indx_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9902 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9910 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9886 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9913 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9891 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9890 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9888 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9889 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9902 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9903 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9884 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add3/U17  ( .Z(\SADR/pgaddxyz[22] ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9904 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9883 ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9887 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9907 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9896 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9899 ), .A(\SADR/pgaddyz[19] ), .B(
        \pk_indx_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9893 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9913 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9897 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9908 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9888 ), .A(\SADR/pgaddyz[23] ), .B(
        \pk_indx_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9895 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9885 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9909 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9901 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9892 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9893 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9886 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add3/U19  ( .Z(\SADR/pgaddxyz[20] ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9906 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9894 ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add3/n9910 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9901 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9887 ), .C(
        \SADR/ADDIDX/add_x_y_z/add3/n9907 ), .D(
        \SADR/ADDIDX/add_x_y_z/add3/n9908 ), .E(
        \SADR/ADDIDX/add_x_y_z/add3/n9911 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9912 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9886 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add3/U16  ( .Z(\SADR/pgaddxyz[23] ), .A(
        \SADR/ADDIDX/add_x_y_z/c_last ), .B(\SADR/ADDIDX/add_x_y_z/add3/n9891 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y_z/add3/U18  ( .Z(\SADR/pgaddxyz[21] ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9905 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9892 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9886 ), .A(\SADR/pgaddyz[21] ), .B(
        \pk_indx_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_x_y_z/add3/n9890 ), .A(\SADR/pgaddyz[23] ), .B(
        \pk_indx_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9908 ), .A(\SADR/pgaddyz[19] ), .B(
        \pk_indx_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9909 ), .A(
        \SADR/ADDIDX/add_x_y_z/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9911 ), .A(\SADR/pgaddyz[20] ), .B(
        \pk_indx_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9913 ), .A(\SADR/pgaddyz[21] ), .B(
        \pk_indx_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y_z/add3/n9904 ), .A(
        \SADR/ADDIDX/add_x_y_z/add3/n9903 ), .B(
        \SADR/ADDIDX/add_x_y_z/add3/n9884 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_z/add0/n9849 ), .B(\SADR/ADDIDX/add_w_z/add0/n9850 
        ), .C(\SADR/ADDIDX/add_w_z/add0/n9851 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_z/add0/n9852 ), .B(\SADR/ADDIDX/add_w_z/add0/n9849 
        ), .C(\SADR/ADDIDX/add_w_z/add0/n9853 ), .D(
        \SADR/ADDIDX/add_w_z/add0/n9854 ), .E(\SADR/ADDIDX/add_w_z/add0/n9855 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9865 ), .A(\SADR/ADDIDX/add_w_z/add0/n9864 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9866 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_z/add0/n9867 ), .A(\SADR/ADDIDX/add_w_z/add0/n9852 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9868 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9868 ), .A(\pk_indw_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9870 ), .A(\SADR/ADDIDX/add_w_z/add0/n9849 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9863 ), .A(\SADR/ADDIDX/add_w_z/add0/n9866 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9852 ), .A(\pk_indw_h[0] ), .B(
        \pk_indz_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9851 ), .A(\pk_indw_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9873 ), .A(\SADR/ADDIDX/add_w_z/add0/n9874 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9878 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add0/U26  ( .Z(\SADR/pgaddwz[0] ), .A(1'b0
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9867 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_z/gg_out[0] ), .A(\SADR/ADDIDX/add_w_z/add0/n9855 ), 
        .B(\SADR/ADDIDX/add_w_z/add0/n9856 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9857 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9861 ), .A(\SADR/ADDIDX/add_w_z/add0/n9862 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9863 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9864 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9872 ), .A(\SADR/ADDIDX/add_w_z/add0/n9876 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9852 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9854 ), .D(\SADR/ADDIDX/add_w_z/add0/n9877 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9849 ), .A(\pk_indw_h[4] ), .B(
        \pk_indz_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9850 ), .A(\SADR/ADDIDX/add_w_z/add0/n9872 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9879 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9860 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add0/U20  ( .Z(\SADR/pgaddwz[1] ), .A(
        \SADR/ADDIDX/add_w_z/add0/n9862 ), .B(\SADR/ADDIDX/add_w_z/add0/n9865 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9874 ), .A(\pk_indw_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9869 ), .A(\SADR/ADDIDX/add_w_z/add0/n9877 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9853 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9880 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9858 ), .A(\SADR/ADDIDX/add_w_z/add0/n9857 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9855 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9856 ), .A(\SADR/ADDIDX/add_w_z/add0/n9869 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9870 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9851 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add0/U17  ( .Z(\SADR/pgaddwz[4] ), .A(
        \SADR/ADDIDX/add_w_z/add0/n9871 ), .B(\SADR/ADDIDX/add_w_z/add0/n9850 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9854 ), .A(\SADR/ADDIDX/add_w_z/add0/n9874 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9863 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9866 ), .A(\pk_indw_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9860 ), .A(\SADR/ADDIDX/add_w_z/add0/n9880 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9864 ), .A(\SADR/ADDIDX/add_w_z/add0/n9875 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9855 ), .A(\pk_indw_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9862 ), .A(\SADR/ADDIDX/add_w_z/add0/n9852 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9876 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9868 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9859 ), .A(\SADR/ADDIDX/add_w_z/add0/n9860 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9853 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add0/U19  ( .Z(\SADR/pgaddwz[2] ), .A(
        \SADR/ADDIDX/add_w_z/add0/n9873 ), .B(\SADR/ADDIDX/add_w_z/add0/n9861 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_z/add0/n9877 ), .A(\SADR/ADDIDX/add_w_z/add0/n9868 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9854 ), .C(
        \SADR/ADDIDX/add_w_z/add0/n9874 ), .D(\SADR/ADDIDX/add_w_z/add0/n9875 
        ), .E(\SADR/ADDIDX/add_w_z/add0/n9878 ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9879 ), .A(\SADR/ADDIDX/add_w_z/add0/n9853 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add0/U16  ( .Z(\SADR/pgaddwz[5] ), .A(
        \SADR/ADDIDX/add_w_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_z/add0/n9858 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add0/U18  ( .Z(\SADR/pgaddwz[3] ), .A(
        \SADR/ADDIDX/add_w_z/add0/n9872 ), .B(\SADR/ADDIDX/add_w_z/add0/n9859 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9853 ), .A(\pk_indw_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_z/add0/n9857 ), .A(\pk_indw_h[5] ), .B(
        \pk_indz_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9875 ), .A(\pk_indw_h[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9876 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9878 ), .A(\pk_indw_h[2] ), .B(
        \pk_indz_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9880 ), .A(\pk_indw_h[3] ), .B(
        \pk_indz_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_z/add0/n9871 ), .A(\SADR/ADDIDX/add_w_z/add0/n9870 
        ), .B(\SADR/ADDIDX/add_w_z/add0/n9851 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_z/add1/n9817 ), .B(\SADR/ADDIDX/add_w_z/add1/n9818 
        ), .C(\SADR/ADDIDX/add_w_z/add1/n9819 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_z/gp_out[1] ), .A(\SADR/ADDIDX/add_w_z/add1/n9820 ), 
        .B(\SADR/ADDIDX/add_w_z/add1/n9817 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9821 ), .D(\SADR/ADDIDX/add_w_z/add1/n9822 
        ), .E(\SADR/ADDIDX/add_w_z/add1/n9823 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9833 ), .A(\SADR/ADDIDX/add_w_z/add1/n9832 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9834 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_z/add1/n9835 ), .A(\SADR/ADDIDX/add_w_z/add1/n9820 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9836 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9836 ), .A(\pk_indw_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9838 ), .A(\SADR/ADDIDX/add_w_z/add1/n9817 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9831 ), .A(\SADR/ADDIDX/add_w_z/add1/n9834 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9820 ), .A(\pk_indw_h[6] ), .B(
        \pk_indz_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9819 ), .A(\pk_indw_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9841 ), .A(\SADR/ADDIDX/add_w_z/add1/n9842 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9846 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add1/U26  ( .Z(\SADR/pgaddwz[6] ), .A(
        \SADR/ADDIDX/add_w_z/gg_out[0] ), .B(\SADR/ADDIDX/add_w_z/add1/n9835 )
         );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_z/gg_out[1] ), .A(\SADR/ADDIDX/add_w_z/add1/n9823 ), 
        .B(\SADR/ADDIDX/add_w_z/add1/n9824 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9825 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9829 ), .A(\SADR/ADDIDX/add_w_z/add1/n9830 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9831 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9832 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9840 ), .A(\SADR/ADDIDX/add_w_z/add1/n9844 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9820 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9822 ), .D(\SADR/ADDIDX/add_w_z/add1/n9845 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9817 ), .A(\pk_indw_h[10] ), .B(
        \pk_indz_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9818 ), .A(\SADR/ADDIDX/add_w_z/add1/n9840 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9847 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9828 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add1/U20  ( .Z(\SADR/pgaddwz[7] ), .A(
        \SADR/ADDIDX/add_w_z/add1/n9830 ), .B(\SADR/ADDIDX/add_w_z/add1/n9833 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9842 ), .A(\pk_indw_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9837 ), .A(\SADR/ADDIDX/add_w_z/add1/n9845 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9821 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9848 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9826 ), .A(\SADR/ADDIDX/add_w_z/add1/n9825 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9823 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9824 ), .A(\SADR/ADDIDX/add_w_z/add1/n9837 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9838 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9819 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add1/U17  ( .Z(\SADR/pgaddwz[10] ), .A(
        \SADR/ADDIDX/add_w_z/add1/n9839 ), .B(\SADR/ADDIDX/add_w_z/add1/n9818 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9822 ), .A(\SADR/ADDIDX/add_w_z/add1/n9842 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9831 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9834 ), .A(\pk_indw_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9828 ), .A(\SADR/ADDIDX/add_w_z/add1/n9848 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9832 ), .A(\SADR/ADDIDX/add_w_z/add1/n9843 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9823 ), .A(\pk_indw_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9830 ), .A(\SADR/ADDIDX/add_w_z/add1/n9820 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9844 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9836 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9827 ), .A(\SADR/ADDIDX/add_w_z/add1/n9828 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9821 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add1/U19  ( .Z(\SADR/pgaddwz[8] ), .A(
        \SADR/ADDIDX/add_w_z/add1/n9841 ), .B(\SADR/ADDIDX/add_w_z/add1/n9829 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_z/add1/n9845 ), .A(\SADR/ADDIDX/add_w_z/add1/n9836 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9822 ), .C(
        \SADR/ADDIDX/add_w_z/add1/n9842 ), .D(\SADR/ADDIDX/add_w_z/add1/n9843 
        ), .E(\SADR/ADDIDX/add_w_z/add1/n9846 ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9847 ), .A(\SADR/ADDIDX/add_w_z/add1/n9821 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add1/U16  ( .Z(\SADR/pgaddwz[11] ), .A(
        \SADR/ADDIDX/add_w_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_z/add1/n9826 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add1/U18  ( .Z(\SADR/pgaddwz[9] ), .A(
        \SADR/ADDIDX/add_w_z/add1/n9840 ), .B(\SADR/ADDIDX/add_w_z/add1/n9827 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9821 ), .A(\pk_indw_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_z/add1/n9825 ), .A(\pk_indw_h[11] ), .B(
        \pk_indz_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9843 ), .A(\pk_indw_h[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9844 ), .A(\SADR/ADDIDX/add_w_z/gg_out[0] )
         );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9846 ), .A(\pk_indw_h[8] ), .B(
        \pk_indz_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9848 ), .A(\pk_indw_h[9] ), .B(
        \pk_indz_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_z/add1/n9839 ), .A(\SADR/ADDIDX/add_w_z/add1/n9838 
        ), .B(\SADR/ADDIDX/add_w_z/add1/n9819 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_z/add2/n9785 ), .B(\SADR/ADDIDX/add_w_z/add2/n9786 
        ), .C(\SADR/ADDIDX/add_w_z/add2/n9787 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_z/gp_out[2] ), .A(\SADR/ADDIDX/add_w_z/add2/n9788 ), 
        .B(\SADR/ADDIDX/add_w_z/add2/n9785 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9789 ), .D(\SADR/ADDIDX/add_w_z/add2/n9790 
        ), .E(\SADR/ADDIDX/add_w_z/add2/n9791 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9801 ), .A(\SADR/ADDIDX/add_w_z/add2/n9800 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9802 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_z/add2/n9803 ), .A(\SADR/ADDIDX/add_w_z/add2/n9788 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9804 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9804 ), .A(\pk_indw_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9806 ), .A(\SADR/ADDIDX/add_w_z/add2/n9785 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9799 ), .A(\SADR/ADDIDX/add_w_z/add2/n9802 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9788 ), .A(\pk_indw_h[12] ), .B(
        \pk_indz_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9787 ), .A(\pk_indw_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9809 ), .A(\SADR/ADDIDX/add_w_z/add2/n9810 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9814 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add2/U26  ( .Z(\SADR/pgaddwz[12] ), .A(
        \SADR/ADDIDX/add_w_z/cin_stg[1] ), .B(\SADR/ADDIDX/add_w_z/add2/n9803 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_z/gg_out[2] ), .A(\SADR/ADDIDX/add_w_z/add2/n9791 ), 
        .B(\SADR/ADDIDX/add_w_z/add2/n9792 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9793 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9797 ), .A(\SADR/ADDIDX/add_w_z/add2/n9798 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9799 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9800 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9808 ), .A(\SADR/ADDIDX/add_w_z/add2/n9812 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9788 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9790 ), .D(\SADR/ADDIDX/add_w_z/add2/n9813 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9785 ), .A(\pk_indw_h[16] ), .B(
        \pk_indz_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9786 ), .A(\SADR/ADDIDX/add_w_z/add2/n9808 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9815 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9796 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add2/U20  ( .Z(\SADR/pgaddwz[13] ), .A(
        \SADR/ADDIDX/add_w_z/add2/n9798 ), .B(\SADR/ADDIDX/add_w_z/add2/n9801 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9810 ), .A(\pk_indw_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9805 ), .A(\SADR/ADDIDX/add_w_z/add2/n9813 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9789 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9816 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9794 ), .A(\SADR/ADDIDX/add_w_z/add2/n9793 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9791 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9792 ), .A(\SADR/ADDIDX/add_w_z/add2/n9805 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9806 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9787 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add2/U17  ( .Z(\SADR/pgaddwz[16] ), .A(
        \SADR/ADDIDX/add_w_z/add2/n9807 ), .B(\SADR/ADDIDX/add_w_z/add2/n9786 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9790 ), .A(\SADR/ADDIDX/add_w_z/add2/n9810 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9799 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9802 ), .A(\pk_indw_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9796 ), .A(\SADR/ADDIDX/add_w_z/add2/n9816 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9800 ), .A(\SADR/ADDIDX/add_w_z/add2/n9811 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9791 ), .A(\pk_indw_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9798 ), .A(\SADR/ADDIDX/add_w_z/add2/n9788 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9812 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9804 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9795 ), .A(\SADR/ADDIDX/add_w_z/add2/n9796 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9789 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add2/U19  ( .Z(\SADR/pgaddwz[14] ), .A(
        \SADR/ADDIDX/add_w_z/add2/n9809 ), .B(\SADR/ADDIDX/add_w_z/add2/n9797 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_z/add2/n9813 ), .A(\SADR/ADDIDX/add_w_z/add2/n9804 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9790 ), .C(
        \SADR/ADDIDX/add_w_z/add2/n9810 ), .D(\SADR/ADDIDX/add_w_z/add2/n9811 
        ), .E(\SADR/ADDIDX/add_w_z/add2/n9814 ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9815 ), .A(\SADR/ADDIDX/add_w_z/add2/n9789 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add2/U16  ( .Z(\SADR/pgaddwz[17] ), .A(
        \SADR/ADDIDX/add_w_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_z/add2/n9794 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add2/U18  ( .Z(\SADR/pgaddwz[15] ), .A(
        \SADR/ADDIDX/add_w_z/add2/n9808 ), .B(\SADR/ADDIDX/add_w_z/add2/n9795 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9789 ), .A(\pk_indw_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_z/add2/n9793 ), .A(\pk_indw_h[17] ), .B(
        \pk_indz_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9811 ), .A(\pk_indw_h[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9812 ), .A(\SADR/ADDIDX/add_w_z/cin_stg[1] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9814 ), .A(\pk_indw_h[14] ), .B(
        \pk_indz_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9816 ), .A(\pk_indw_h[15] ), .B(
        \pk_indz_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_z/add2/n9807 ), .A(\SADR/ADDIDX/add_w_z/add2/n9806 
        ), .B(\SADR/ADDIDX/add_w_z/add2/n9787 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_z/c_last ), .A(\SADR/ADDIDX/add_w_z/add3/n9753 ), 
        .B(\SADR/ADDIDX/add_w_z/add3/n9754 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9755 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_z/gp_out[3] ), .A(\SADR/ADDIDX/add_w_z/add3/n9756 ), 
        .B(\SADR/ADDIDX/add_w_z/add3/n9753 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9757 ), .D(\SADR/ADDIDX/add_w_z/add3/n9758 
        ), .E(\SADR/ADDIDX/add_w_z/add3/n9759 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9769 ), .A(\SADR/ADDIDX/add_w_z/add3/n9768 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9770 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_z/add3/n9771 ), .A(\SADR/ADDIDX/add_w_z/add3/n9756 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9772 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9772 ), .A(\pk_indw_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9774 ), .A(\SADR/ADDIDX/add_w_z/add3/n9753 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9767 ), .A(\SADR/ADDIDX/add_w_z/add3/n9770 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9756 ), .A(\pk_indw_h[18] ), .B(
        \pk_indz_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9755 ), .A(\pk_indw_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9777 ), .A(\SADR/ADDIDX/add_w_z/add3/n9778 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9782 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add3/U26  ( .Z(\SADR/pgaddwz[18] ), .A(
        \SADR/ADDIDX/add_w_z/cin_stg[2] ), .B(\SADR/ADDIDX/add_w_z/add3/n9771 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_z/gg_out[3] ), .A(\SADR/ADDIDX/add_w_z/add3/n9759 ), 
        .B(\SADR/ADDIDX/add_w_z/add3/n9760 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9761 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9765 ), .A(\SADR/ADDIDX/add_w_z/add3/n9766 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9767 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9768 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9776 ), .A(\SADR/ADDIDX/add_w_z/add3/n9780 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9756 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9758 ), .D(\SADR/ADDIDX/add_w_z/add3/n9781 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9753 ), .A(\pk_indw_h[22] ), .B(
        \pk_indz_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9754 ), .A(\SADR/ADDIDX/add_w_z/add3/n9776 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9783 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9764 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add3/U20  ( .Z(\SADR/pgaddwz[19] ), .A(
        \SADR/ADDIDX/add_w_z/add3/n9766 ), .B(\SADR/ADDIDX/add_w_z/add3/n9769 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9778 ), .A(\pk_indw_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9773 ), .A(\SADR/ADDIDX/add_w_z/add3/n9781 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9757 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9784 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9762 ), .A(\SADR/ADDIDX/add_w_z/add3/n9761 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9759 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9760 ), .A(\SADR/ADDIDX/add_w_z/add3/n9773 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9774 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9755 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add3/U17  ( .Z(\SADR/pgaddwz[22] ), .A(
        \SADR/ADDIDX/add_w_z/add3/n9775 ), .B(\SADR/ADDIDX/add_w_z/add3/n9754 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9758 ), .A(\SADR/ADDIDX/add_w_z/add3/n9778 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9767 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9770 ), .A(\pk_indw_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9764 ), .A(\SADR/ADDIDX/add_w_z/add3/n9784 
        ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9768 ), .A(\SADR/ADDIDX/add_w_z/add3/n9779 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9759 ), .A(\pk_indw_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9766 ), .A(\SADR/ADDIDX/add_w_z/add3/n9756 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9780 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9772 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9763 ), .A(\SADR/ADDIDX/add_w_z/add3/n9764 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9757 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add3/U19  ( .Z(\SADR/pgaddwz[20] ), .A(
        \SADR/ADDIDX/add_w_z/add3/n9777 ), .B(\SADR/ADDIDX/add_w_z/add3/n9765 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_z/add3/n9781 ), .A(\SADR/ADDIDX/add_w_z/add3/n9772 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9758 ), .C(
        \SADR/ADDIDX/add_w_z/add3/n9778 ), .D(\SADR/ADDIDX/add_w_z/add3/n9779 
        ), .E(\SADR/ADDIDX/add_w_z/add3/n9782 ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9783 ), .A(\SADR/ADDIDX/add_w_z/add3/n9757 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add3/U16  ( .Z(\SADR/pgaddwz[23] ), .A(
        \SADR/ADDIDX/add_w_z/c_last ), .B(\SADR/ADDIDX/add_w_z/add3/n9762 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_z/add3/U18  ( .Z(\SADR/pgaddwz[21] ), .A(
        \SADR/ADDIDX/add_w_z/add3/n9776 ), .B(\SADR/ADDIDX/add_w_z/add3/n9763 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9757 ), .A(\pk_indw_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_z/add3/n9761 ), .A(\pk_indw_h[23] ), .B(
        \pk_indz_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9779 ), .A(\pk_indw_h[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9780 ), .A(\SADR/ADDIDX/add_w_z/cin_stg[2] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9782 ), .A(\pk_indw_h[20] ), .B(
        \pk_indz_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9784 ), .A(\pk_indw_h[21] ), .B(
        \pk_indz_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_z/add3/n9775 ), .A(\SADR/ADDIDX/add_w_z/add3/n9774 
        ), .B(\SADR/ADDIDX/add_w_z/add3/n9755 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/c_last ), .A(
        \SADR/ADDIDX/add_x_y/add0/n9720 ), .B(\SADR/ADDIDX/add_x_y/add0/n9721 
        ), .C(\SADR/ADDIDX/add_x_y/add0/n9722 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/gp_out ), .A(
        \SADR/ADDIDX/add_x_y/add0/n9723 ), .B(\SADR/ADDIDX/add_x_y/add0/n9720 
        ), .C(\SADR/ADDIDX/add_x_y/add0/n9724 ), .D(
        \SADR/ADDIDX/add_x_y/add0/n9725 ), .E(\SADR/ADDIDX/add_x_y/add0/n9726 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9736 ), .A(\SADR/ADDIDX/add_x_y/add0/n9735 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9737 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y/add0/U14  ( .Z(
        \SADR/ADDIDX/add_x_y/add0/n9738 ), .A(\SADR/ADDIDX/add_x_y/add0/n9723 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9739 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9739 ), .A(\pk_indx_h[0] ), .B(
        \pk_indy_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9741 ), .A(\SADR/ADDIDX/add_x_y/add0/n9720 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9734 ), .A(\SADR/ADDIDX/add_x_y/add0/n9737 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9723 ), .A(\pk_indx_h[0] ), .B(
        \pk_indy_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9722 ), .A(\pk_indx_h[4] ), .B(
        \pk_indy_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9744 ), .A(\SADR/ADDIDX/add_x_y/add0/n9745 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9749 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add0/U26  ( .Z(\SADR/pgaddxy[0] ), .A(1'b0
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9738 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y/add0/U9  ( .Z(
        \SADR/ADDIDX/add_x_y/gg_out[0] ), .A(\SADR/ADDIDX/add_x_y/add0/n9726 ), 
        .B(\SADR/ADDIDX/add_x_y/add0/n9727 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9728 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9732 ), .A(\SADR/ADDIDX/add_x_y/add0/n9733 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9734 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9735 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9743 ), .A(\SADR/ADDIDX/add_x_y/add0/n9747 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9723 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9725 ), .D(\SADR/ADDIDX/add_x_y/add0/n9748 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9720 ), .A(\pk_indx_h[4] ), .B(
        \pk_indy_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9721 ), .A(\SADR/ADDIDX/add_x_y/add0/n9743 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9750 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9731 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add0/U20  ( .Z(\SADR/pgaddxy[1] ), .A(
        \SADR/ADDIDX/add_x_y/add0/n9733 ), .B(\SADR/ADDIDX/add_x_y/add0/n9736 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9745 ), .A(\pk_indx_h[2] ), .B(
        \pk_indy_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9740 ), .A(\SADR/ADDIDX/add_x_y/add0/n9748 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9724 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9751 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9729 ), .A(\SADR/ADDIDX/add_x_y/add0/n9728 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9726 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9727 ), .A(\SADR/ADDIDX/add_x_y/add0/n9740 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9741 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9722 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add0/U17  ( .Z(\SADR/pgaddxy[4] ), .A(
        \SADR/ADDIDX/add_x_y/add0/n9742 ), .B(\SADR/ADDIDX/add_x_y/add0/n9721 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9725 ), .A(\SADR/ADDIDX/add_x_y/add0/n9745 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9734 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9737 ), .A(\pk_indx_h[1] ), .B(
        \pk_indy_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9731 ), .A(\SADR/ADDIDX/add_x_y/add0/n9751 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9735 ), .A(\SADR/ADDIDX/add_x_y/add0/n9746 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9726 ), .A(\pk_indx_h[5] ), .B(
        \pk_indy_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9733 ), .A(\SADR/ADDIDX/add_x_y/add0/n9723 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9747 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9739 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9730 ), .A(\SADR/ADDIDX/add_x_y/add0/n9731 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9724 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add0/U19  ( .Z(\SADR/pgaddxy[2] ), .A(
        \SADR/ADDIDX/add_x_y/add0/n9744 ), .B(\SADR/ADDIDX/add_x_y/add0/n9732 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y/add0/U25  ( .Z(
        \SADR/ADDIDX/add_x_y/add0/n9748 ), .A(\SADR/ADDIDX/add_x_y/add0/n9739 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9725 ), .C(
        \SADR/ADDIDX/add_x_y/add0/n9745 ), .D(\SADR/ADDIDX/add_x_y/add0/n9746 
        ), .E(\SADR/ADDIDX/add_x_y/add0/n9749 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9750 ), .A(\SADR/ADDIDX/add_x_y/add0/n9724 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add0/U16  ( .Z(\SADR/pgaddxy[5] ), .A(
        \SADR/ADDIDX/add_x_y/add0/c_last ), .B(
        \SADR/ADDIDX/add_x_y/add0/n9729 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add0/U18  ( .Z(\SADR/pgaddxy[3] ), .A(
        \SADR/ADDIDX/add_x_y/add0/n9743 ), .B(\SADR/ADDIDX/add_x_y/add0/n9730 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9724 ), .A(\pk_indx_h[3] ), .B(
        \pk_indy_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y/add0/U43  ( .Z(
        \SADR/ADDIDX/add_x_y/add0/n9728 ), .A(\pk_indx_h[5] ), .B(
        \pk_indy_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9746 ), .A(\pk_indx_h[1] ), .B(
        \pk_indy_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9747 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9749 ), .A(\pk_indx_h[2] ), .B(
        \pk_indy_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9751 ), .A(\pk_indx_h[3] ), .B(
        \pk_indy_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y/add0/n9742 ), .A(\SADR/ADDIDX/add_x_y/add0/n9741 
        ), .B(\SADR/ADDIDX/add_x_y/add0/n9722 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/c_last ), .A(
        \SADR/ADDIDX/add_x_y/add1/n9688 ), .B(\SADR/ADDIDX/add_x_y/add1/n9689 
        ), .C(\SADR/ADDIDX/add_x_y/add1/n9690 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y/gp_out[1] ), .A(\SADR/ADDIDX/add_x_y/add1/n9691 ), 
        .B(\SADR/ADDIDX/add_x_y/add1/n9688 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9692 ), .D(\SADR/ADDIDX/add_x_y/add1/n9693 
        ), .E(\SADR/ADDIDX/add_x_y/add1/n9694 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9704 ), .A(\SADR/ADDIDX/add_x_y/add1/n9703 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9705 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y/add1/U14  ( .Z(
        \SADR/ADDIDX/add_x_y/add1/n9706 ), .A(\SADR/ADDIDX/add_x_y/add1/n9691 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9707 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9707 ), .A(\pk_indx_h[6] ), .B(
        \pk_indy_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9709 ), .A(\SADR/ADDIDX/add_x_y/add1/n9688 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9702 ), .A(\SADR/ADDIDX/add_x_y/add1/n9705 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9691 ), .A(\pk_indx_h[6] ), .B(
        \pk_indy_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9690 ), .A(\pk_indx_h[10] ), .B(
        \pk_indy_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9712 ), .A(\SADR/ADDIDX/add_x_y/add1/n9713 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9717 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add1/U26  ( .Z(\SADR/pgaddxy[6] ), .A(
        \SADR/ADDIDX/add_x_y/gg_out[0] ), .B(\SADR/ADDIDX/add_x_y/add1/n9706 )
         );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y/add1/U9  ( .Z(
        \SADR/ADDIDX/add_x_y/gg_out[1] ), .A(\SADR/ADDIDX/add_x_y/add1/n9694 ), 
        .B(\SADR/ADDIDX/add_x_y/add1/n9695 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9696 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9700 ), .A(\SADR/ADDIDX/add_x_y/add1/n9701 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9702 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9703 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9711 ), .A(\SADR/ADDIDX/add_x_y/add1/n9715 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9691 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9693 ), .D(\SADR/ADDIDX/add_x_y/add1/n9716 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9688 ), .A(\pk_indx_h[10] ), .B(
        \pk_indy_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9689 ), .A(\SADR/ADDIDX/add_x_y/add1/n9711 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9718 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9699 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add1/U20  ( .Z(\SADR/pgaddxy[7] ), .A(
        \SADR/ADDIDX/add_x_y/add1/n9701 ), .B(\SADR/ADDIDX/add_x_y/add1/n9704 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9713 ), .A(\pk_indx_h[8] ), .B(
        \pk_indy_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9708 ), .A(\SADR/ADDIDX/add_x_y/add1/n9716 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9692 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9719 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9697 ), .A(\SADR/ADDIDX/add_x_y/add1/n9696 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9694 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9695 ), .A(\SADR/ADDIDX/add_x_y/add1/n9708 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9709 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9690 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add1/U17  ( .Z(\SADR/pgaddxy[10] ), .A(
        \SADR/ADDIDX/add_x_y/add1/n9710 ), .B(\SADR/ADDIDX/add_x_y/add1/n9689 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9693 ), .A(\SADR/ADDIDX/add_x_y/add1/n9713 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9702 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9705 ), .A(\pk_indx_h[7] ), .B(
        \pk_indy_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9699 ), .A(\SADR/ADDIDX/add_x_y/add1/n9719 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9703 ), .A(\SADR/ADDIDX/add_x_y/add1/n9714 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9694 ), .A(\pk_indx_h[11] ), .B(
        \pk_indy_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9701 ), .A(\SADR/ADDIDX/add_x_y/add1/n9691 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9715 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9707 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9698 ), .A(\SADR/ADDIDX/add_x_y/add1/n9699 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9692 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add1/U19  ( .Z(\SADR/pgaddxy[8] ), .A(
        \SADR/ADDIDX/add_x_y/add1/n9712 ), .B(\SADR/ADDIDX/add_x_y/add1/n9700 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y/add1/U25  ( .Z(
        \SADR/ADDIDX/add_x_y/add1/n9716 ), .A(\SADR/ADDIDX/add_x_y/add1/n9707 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9693 ), .C(
        \SADR/ADDIDX/add_x_y/add1/n9713 ), .D(\SADR/ADDIDX/add_x_y/add1/n9714 
        ), .E(\SADR/ADDIDX/add_x_y/add1/n9717 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9718 ), .A(\SADR/ADDIDX/add_x_y/add1/n9692 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add1/U16  ( .Z(\SADR/pgaddxy[11] ), .A(
        \SADR/ADDIDX/add_x_y/add1/c_last ), .B(
        \SADR/ADDIDX/add_x_y/add1/n9697 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add1/U18  ( .Z(\SADR/pgaddxy[9] ), .A(
        \SADR/ADDIDX/add_x_y/add1/n9711 ), .B(\SADR/ADDIDX/add_x_y/add1/n9698 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9692 ), .A(\pk_indx_h[9] ), .B(
        \pk_indy_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y/add1/U43  ( .Z(
        \SADR/ADDIDX/add_x_y/add1/n9696 ), .A(\pk_indx_h[11] ), .B(
        \pk_indy_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9714 ), .A(\pk_indx_h[7] ), .B(
        \pk_indy_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9715 ), .A(\SADR/ADDIDX/add_x_y/gg_out[0] )
         );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9717 ), .A(\pk_indx_h[8] ), .B(
        \pk_indy_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9719 ), .A(\pk_indx_h[9] ), .B(
        \pk_indy_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y/add1/n9710 ), .A(\SADR/ADDIDX/add_x_y/add1/n9709 
        ), .B(\SADR/ADDIDX/add_x_y/add1/n9690 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/c_last ), .A(
        \SADR/ADDIDX/add_x_y/add2/n9656 ), .B(\SADR/ADDIDX/add_x_y/add2/n9657 
        ), .C(\SADR/ADDIDX/add_x_y/add2/n9658 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y/gp_out[2] ), .A(\SADR/ADDIDX/add_x_y/add2/n9659 ), 
        .B(\SADR/ADDIDX/add_x_y/add2/n9656 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9660 ), .D(\SADR/ADDIDX/add_x_y/add2/n9661 
        ), .E(\SADR/ADDIDX/add_x_y/add2/n9662 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9672 ), .A(\SADR/ADDIDX/add_x_y/add2/n9671 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9673 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y/add2/U14  ( .Z(
        \SADR/ADDIDX/add_x_y/add2/n9674 ), .A(\SADR/ADDIDX/add_x_y/add2/n9659 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9675 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9675 ), .A(\pk_indx_h[12] ), .B(
        \pk_indy_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9677 ), .A(\SADR/ADDIDX/add_x_y/add2/n9656 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9670 ), .A(\SADR/ADDIDX/add_x_y/add2/n9673 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9659 ), .A(\pk_indx_h[12] ), .B(
        \pk_indy_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9658 ), .A(\pk_indx_h[16] ), .B(
        \pk_indy_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9680 ), .A(\SADR/ADDIDX/add_x_y/add2/n9681 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9685 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add2/U26  ( .Z(\SADR/pgaddxy[12] ), .A(
        \SADR/ADDIDX/add_x_y/cin_stg[1] ), .B(\SADR/ADDIDX/add_x_y/add2/n9674 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y/add2/U9  ( .Z(
        \SADR/ADDIDX/add_x_y/gg_out[2] ), .A(\SADR/ADDIDX/add_x_y/add2/n9662 ), 
        .B(\SADR/ADDIDX/add_x_y/add2/n9663 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9664 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9668 ), .A(\SADR/ADDIDX/add_x_y/add2/n9669 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9670 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9671 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9679 ), .A(\SADR/ADDIDX/add_x_y/add2/n9683 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9659 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9661 ), .D(\SADR/ADDIDX/add_x_y/add2/n9684 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9656 ), .A(\pk_indx_h[16] ), .B(
        \pk_indy_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9657 ), .A(\SADR/ADDIDX/add_x_y/add2/n9679 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9686 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9667 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add2/U20  ( .Z(\SADR/pgaddxy[13] ), .A(
        \SADR/ADDIDX/add_x_y/add2/n9669 ), .B(\SADR/ADDIDX/add_x_y/add2/n9672 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9681 ), .A(\pk_indx_h[14] ), .B(
        \pk_indy_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9676 ), .A(\SADR/ADDIDX/add_x_y/add2/n9684 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9660 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9687 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9665 ), .A(\SADR/ADDIDX/add_x_y/add2/n9664 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9662 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9663 ), .A(\SADR/ADDIDX/add_x_y/add2/n9676 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9677 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9658 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add2/U17  ( .Z(\SADR/pgaddxy[16] ), .A(
        \SADR/ADDIDX/add_x_y/add2/n9678 ), .B(\SADR/ADDIDX/add_x_y/add2/n9657 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9661 ), .A(\SADR/ADDIDX/add_x_y/add2/n9681 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9670 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9673 ), .A(\pk_indx_h[13] ), .B(
        \pk_indy_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9667 ), .A(\SADR/ADDIDX/add_x_y/add2/n9687 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9671 ), .A(\SADR/ADDIDX/add_x_y/add2/n9682 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9662 ), .A(\pk_indx_h[17] ), .B(
        \pk_indy_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9669 ), .A(\SADR/ADDIDX/add_x_y/add2/n9659 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9683 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9675 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9666 ), .A(\SADR/ADDIDX/add_x_y/add2/n9667 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9660 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add2/U19  ( .Z(\SADR/pgaddxy[14] ), .A(
        \SADR/ADDIDX/add_x_y/add2/n9680 ), .B(\SADR/ADDIDX/add_x_y/add2/n9668 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y/add2/U25  ( .Z(
        \SADR/ADDIDX/add_x_y/add2/n9684 ), .A(\SADR/ADDIDX/add_x_y/add2/n9675 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9661 ), .C(
        \SADR/ADDIDX/add_x_y/add2/n9681 ), .D(\SADR/ADDIDX/add_x_y/add2/n9682 
        ), .E(\SADR/ADDIDX/add_x_y/add2/n9685 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9686 ), .A(\SADR/ADDIDX/add_x_y/add2/n9660 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add2/U16  ( .Z(\SADR/pgaddxy[17] ), .A(
        \SADR/ADDIDX/add_x_y/add2/c_last ), .B(
        \SADR/ADDIDX/add_x_y/add2/n9665 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add2/U18  ( .Z(\SADR/pgaddxy[15] ), .A(
        \SADR/ADDIDX/add_x_y/add2/n9679 ), .B(\SADR/ADDIDX/add_x_y/add2/n9666 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9660 ), .A(\pk_indx_h[15] ), .B(
        \pk_indy_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y/add2/U43  ( .Z(
        \SADR/ADDIDX/add_x_y/add2/n9664 ), .A(\pk_indx_h[17] ), .B(
        \pk_indy_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9682 ), .A(\pk_indx_h[13] ), .B(
        \pk_indy_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9683 ), .A(\SADR/ADDIDX/add_x_y/cin_stg[1] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9685 ), .A(\pk_indx_h[14] ), .B(
        \pk_indy_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9687 ), .A(\pk_indx_h[15] ), .B(
        \pk_indy_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y/add2/n9678 ), .A(\SADR/ADDIDX/add_x_y/add2/n9677 
        ), .B(\SADR/ADDIDX/add_x_y/add2/n9658 ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_x_y/c_last ), .A(\SADR/ADDIDX/add_x_y/add3/n9624 ), 
        .B(\SADR/ADDIDX/add_x_y/add3/n9625 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9626 ) );
    snl_nor05x1 \SADR/ADDIDX/add_x_y/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_x_y/gp_out[3] ), .A(\SADR/ADDIDX/add_x_y/add3/n9627 ), 
        .B(\SADR/ADDIDX/add_x_y/add3/n9624 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9628 ), .D(\SADR/ADDIDX/add_x_y/add3/n9629 
        ), .E(\SADR/ADDIDX/add_x_y/add3/n9630 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9640 ), .A(\SADR/ADDIDX/add_x_y/add3/n9639 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9641 ) );
    snl_and12x1 \SADR/ADDIDX/add_x_y/add3/U14  ( .Z(
        \SADR/ADDIDX/add_x_y/add3/n9642 ), .A(\SADR/ADDIDX/add_x_y/add3/n9627 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9643 ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9643 ), .A(\pk_indx_h[18] ), .B(
        \pk_indy_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9645 ), .A(\SADR/ADDIDX/add_x_y/add3/n9624 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9638 ), .A(\SADR/ADDIDX/add_x_y/add3/n9641 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9627 ), .A(\pk_indx_h[18] ), .B(
        \pk_indy_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9626 ), .A(\pk_indx_h[22] ), .B(
        \pk_indy_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9648 ), .A(\SADR/ADDIDX/add_x_y/add3/n9649 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9653 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add3/U26  ( .Z(\SADR/pgaddxy[18] ), .A(
        \SADR/ADDIDX/add_x_y/cin_stg[2] ), .B(\SADR/ADDIDX/add_x_y/add3/n9642 
        ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_x_y/add3/U9  ( .Z(
        \SADR/ADDIDX/add_x_y/gg_out[3] ), .A(\SADR/ADDIDX/add_x_y/add3/n9630 ), 
        .B(\SADR/ADDIDX/add_x_y/add3/n9631 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9632 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9636 ), .A(\SADR/ADDIDX/add_x_y/add3/n9637 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9638 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9639 ) );
    snl_oai013x0 \SADR/ADDIDX/add_x_y/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9647 ), .A(\SADR/ADDIDX/add_x_y/add3/n9651 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9627 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9629 ), .D(\SADR/ADDIDX/add_x_y/add3/n9652 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9624 ), .A(\pk_indx_h[22] ), .B(
        \pk_indy_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_x_y/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9625 ), .A(\SADR/ADDIDX/add_x_y/add3/n9647 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9654 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9635 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add3/U20  ( .Z(\SADR/pgaddxy[19] ), .A(
        \SADR/ADDIDX/add_x_y/add3/n9637 ), .B(\SADR/ADDIDX/add_x_y/add3/n9640 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9649 ), .A(\pk_indx_h[20] ), .B(
        \pk_indy_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9644 ), .A(\SADR/ADDIDX/add_x_y/add3/n9652 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9628 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9655 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9633 ), .A(\SADR/ADDIDX/add_x_y/add3/n9632 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9630 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_x_y/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9631 ), .A(\SADR/ADDIDX/add_x_y/add3/n9644 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9645 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9626 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add3/U17  ( .Z(\SADR/pgaddxy[22] ), .A(
        \SADR/ADDIDX/add_x_y/add3/n9646 ), .B(\SADR/ADDIDX/add_x_y/add3/n9625 
        ) );
    snl_nand12x1 \SADR/ADDIDX/add_x_y/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9629 ), .A(\SADR/ADDIDX/add_x_y/add3/n9649 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9638 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9641 ), .A(\pk_indx_h[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9635 ), .A(\SADR/ADDIDX/add_x_y/add3/n9655 
        ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9639 ), .A(\SADR/ADDIDX/add_x_y/add3/n9650 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9630 ), .A(\pk_indx_h[23] ), .B(
        \pk_indy_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_x_y/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9637 ), .A(\SADR/ADDIDX/add_x_y/add3/n9627 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9651 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9643 ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9634 ), .A(\SADR/ADDIDX/add_x_y/add3/n9635 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9628 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add3/U19  ( .Z(\SADR/pgaddxy[20] ), .A(
        \SADR/ADDIDX/add_x_y/add3/n9648 ), .B(\SADR/ADDIDX/add_x_y/add3/n9636 
        ) );
    snl_oa122x1 \SADR/ADDIDX/add_x_y/add3/U25  ( .Z(
        \SADR/ADDIDX/add_x_y/add3/n9652 ), .A(\SADR/ADDIDX/add_x_y/add3/n9643 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9629 ), .C(
        \SADR/ADDIDX/add_x_y/add3/n9649 ), .D(\SADR/ADDIDX/add_x_y/add3/n9650 
        ), .E(\SADR/ADDIDX/add_x_y/add3/n9653 ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9654 ), .A(\SADR/ADDIDX/add_x_y/add3/n9628 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add3/U16  ( .Z(\SADR/pgaddxy[23] ), .A(
        \SADR/ADDIDX/add_x_y/c_last ), .B(\SADR/ADDIDX/add_x_y/add3/n9633 ) );
    snl_xor2x0 \SADR/ADDIDX/add_x_y/add3/U18  ( .Z(\SADR/pgaddxy[21] ), .A(
        \SADR/ADDIDX/add_x_y/add3/n9647 ), .B(\SADR/ADDIDX/add_x_y/add3/n9634 
        ) );
    snl_nor02x1 \SADR/ADDIDX/add_x_y/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9628 ), .A(\pk_indx_h[21] ), .B(
        \pk_indy_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_x_y/add3/U43  ( .Z(
        \SADR/ADDIDX/add_x_y/add3/n9632 ), .A(\pk_indx_h[23] ), .B(
        \pk_indy_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9650 ), .A(\pk_indx_h[19] ), .B(
        \pk_indy_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_x_y/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9651 ), .A(\SADR/ADDIDX/add_x_y/cin_stg[2] 
        ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9653 ), .A(\pk_indx_h[20] ), .B(
        \pk_indy_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9655 ), .A(\pk_indx_h[21] ), .B(
        \pk_indy_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_x_y/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_x_y/add3/n9646 ), .A(\SADR/ADDIDX/add_x_y/add3/n9645 
        ), .B(\SADR/ADDIDX/add_x_y/add3/n9626 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9591 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9592 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9593 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9594 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9591 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9595 ), .D(
        \SADR/ADDIDX/add_w_x_z/add0/n9596 ), .E(
        \SADR/ADDIDX/add_w_x_z/add0/n9597 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9607 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9606 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9608 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add0/n9609 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9594 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9610 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9610 ), .A(\SADR/pgaddxz[0] ), .B(
        \pk_indw_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9612 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9591 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9605 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9608 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9594 ), .A(\SADR/pgaddxz[0] ), .B(
        \pk_indw_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9593 ), .A(\SADR/pgaddxz[4] ), .B(
        \pk_indw_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9615 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9616 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9620 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add0/U26  ( .Z(\SADR/pgaddwxz[0] ), .A(
        1'b0), .B(\SADR/ADDIDX/add_w_x_z/add0/n9609 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_z/gg_out[0] ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9597 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9598 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9599 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9603 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9604 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9605 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9606 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9614 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9618 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9594 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9596 ), .D(
        \SADR/ADDIDX/add_w_x_z/add0/n9619 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9591 ), .A(\SADR/pgaddxz[4] ), .B(
        \pk_indw_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9592 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9614 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9621 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9602 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add0/U20  ( .Z(\SADR/pgaddwxz[1] ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9604 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9607 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9616 ), .A(\SADR/pgaddxz[2] ), .B(
        \pk_indw_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9611 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9619 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9595 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9622 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9600 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9599 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9597 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9598 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9611 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9612 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9593 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add0/U17  ( .Z(\SADR/pgaddwxz[4] ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9613 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9592 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9596 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9616 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9605 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9608 ), .A(\SADR/pgaddxz[1] ), .B(
        \pk_indw_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9602 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9622 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9606 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9617 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9597 ), .A(\SADR/pgaddxz[5] ), .B(
        \pk_indw_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9604 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9594 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9618 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9610 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9601 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9602 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9595 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add0/U19  ( .Z(\SADR/pgaddwxz[2] ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9615 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9603 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add0/n9619 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9610 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9596 ), .C(
        \SADR/ADDIDX/add_w_x_z/add0/n9616 ), .D(
        \SADR/ADDIDX/add_w_x_z/add0/n9617 ), .E(
        \SADR/ADDIDX/add_w_x_z/add0/n9620 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9621 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9595 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add0/U16  ( .Z(\SADR/pgaddwxz[5] ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9600 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add0/U18  ( .Z(\SADR/pgaddwxz[3] ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9614 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9601 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9595 ), .A(\SADR/pgaddxz[3] ), .B(
        \pk_indw_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add0/n9599 ), .A(\SADR/pgaddxz[5] ), .B(
        \pk_indw_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9617 ), .A(\SADR/pgaddxz[1] ), .B(
        \pk_indw_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9618 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9620 ), .A(\SADR/pgaddxz[2] ), .B(
        \pk_indw_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9622 ), .A(\SADR/pgaddxz[3] ), .B(
        \pk_indw_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add0/n9613 ), .A(
        \SADR/ADDIDX/add_w_x_z/add0/n9612 ), .B(
        \SADR/ADDIDX/add_w_x_z/add0/n9593 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9559 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9560 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9561 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/gp_out[1] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9562 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9559 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9563 ), .D(
        \SADR/ADDIDX/add_w_x_z/add1/n9564 ), .E(
        \SADR/ADDIDX/add_w_x_z/add1/n9565 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9575 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9574 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9576 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add1/n9577 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9562 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9578 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9578 ), .A(\SADR/pgaddxz[6] ), .B(
        \pk_indw_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9580 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9559 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9573 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9576 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9562 ), .A(\SADR/pgaddxz[6] ), .B(
        \pk_indw_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9561 ), .A(\SADR/pgaddxz[10] ), .B(
        \pk_indw_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9583 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9584 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9588 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add1/U26  ( .Z(\SADR/pgaddwxz[6] ), .A(
        \SADR/ADDIDX/add_w_x_z/gg_out[0] ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9577 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_z/gg_out[1] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9565 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9566 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9567 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9571 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9572 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9573 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9574 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9582 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9586 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9562 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9564 ), .D(
        \SADR/ADDIDX/add_w_x_z/add1/n9587 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9559 ), .A(\SADR/pgaddxz[10] ), .B(
        \pk_indw_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9560 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9582 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9589 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9570 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add1/U20  ( .Z(\SADR/pgaddwxz[7] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9572 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9575 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9584 ), .A(\SADR/pgaddxz[8] ), .B(
        \pk_indw_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9579 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9587 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9563 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9590 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9568 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9567 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9565 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9566 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9579 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9580 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9561 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add1/U17  ( .Z(\SADR/pgaddwxz[10] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9581 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9560 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9564 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9584 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9573 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9576 ), .A(\SADR/pgaddxz[7] ), .B(
        \pk_indw_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9570 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9590 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9574 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9585 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9565 ), .A(\SADR/pgaddxz[11] ), .B(
        \pk_indw_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9572 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9562 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9586 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9578 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9569 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9570 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9563 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add1/U19  ( .Z(\SADR/pgaddwxz[8] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9583 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9571 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add1/n9587 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9578 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9564 ), .C(
        \SADR/ADDIDX/add_w_x_z/add1/n9584 ), .D(
        \SADR/ADDIDX/add_w_x_z/add1/n9585 ), .E(
        \SADR/ADDIDX/add_w_x_z/add1/n9588 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9589 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9563 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add1/U16  ( .Z(\SADR/pgaddwxz[11] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9568 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add1/U18  ( .Z(\SADR/pgaddwxz[9] ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9582 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9569 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9563 ), .A(\SADR/pgaddxz[9] ), .B(
        \pk_indw_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add1/n9567 ), .A(\SADR/pgaddxz[11] ), .B(
        \pk_indw_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9585 ), .A(\SADR/pgaddxz[7] ), .B(
        \pk_indw_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9586 ), .A(
        \SADR/ADDIDX/add_w_x_z/gg_out[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9588 ), .A(\SADR/pgaddxz[8] ), .B(
        \pk_indw_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9590 ), .A(\SADR/pgaddxz[9] ), .B(
        \pk_indw_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add1/n9581 ), .A(
        \SADR/ADDIDX/add_w_x_z/add1/n9580 ), .B(
        \SADR/ADDIDX/add_w_x_z/add1/n9561 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9527 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9528 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9529 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/gp_out[2] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9530 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9527 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9531 ), .D(
        \SADR/ADDIDX/add_w_x_z/add2/n9532 ), .E(
        \SADR/ADDIDX/add_w_x_z/add2/n9533 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9543 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9542 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9544 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add2/n9545 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9530 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9546 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9546 ), .A(\SADR/pgaddxz[12] ), .B(
        \pk_indw_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9548 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9527 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9541 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9544 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9530 ), .A(\SADR/pgaddxz[12] ), .B(
        \pk_indw_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9529 ), .A(\SADR/pgaddxz[16] ), .B(
        \pk_indw_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9551 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9552 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9556 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add2/U26  ( .Z(\SADR/pgaddwxz[12] ), .A(
        \SADR/ADDIDX/add_w_x_z/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9545 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_z/gg_out[2] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9533 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9534 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9535 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9539 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9540 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9541 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9542 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9550 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9554 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9530 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9532 ), .D(
        \SADR/ADDIDX/add_w_x_z/add2/n9555 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9527 ), .A(\SADR/pgaddxz[16] ), .B(
        \pk_indw_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9528 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9550 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9557 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9538 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add2/U20  ( .Z(\SADR/pgaddwxz[13] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9540 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9543 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9552 ), .A(\SADR/pgaddxz[14] ), .B(
        \pk_indw_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9547 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9555 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9531 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9558 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9536 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9535 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9533 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9534 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9547 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9548 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9529 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add2/U17  ( .Z(\SADR/pgaddwxz[16] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9549 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9528 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9532 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9552 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9541 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9544 ), .A(\SADR/pgaddxz[13] ), .B(
        \pk_indw_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9538 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9558 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9542 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9553 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9533 ), .A(\SADR/pgaddxz[17] ), .B(
        \pk_indw_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9540 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9530 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9554 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9546 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9537 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9538 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9531 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add2/U19  ( .Z(\SADR/pgaddwxz[14] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9551 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9539 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add2/n9555 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9546 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9532 ), .C(
        \SADR/ADDIDX/add_w_x_z/add2/n9552 ), .D(
        \SADR/ADDIDX/add_w_x_z/add2/n9553 ), .E(
        \SADR/ADDIDX/add_w_x_z/add2/n9556 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9557 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9531 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add2/U16  ( .Z(\SADR/pgaddwxz[17] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9536 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add2/U18  ( .Z(\SADR/pgaddwxz[15] ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9550 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9537 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9531 ), .A(\SADR/pgaddxz[15] ), .B(
        \pk_indw_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add2/n9535 ), .A(\SADR/pgaddxz[17] ), .B(
        \pk_indw_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9553 ), .A(\SADR/pgaddxz[13] ), .B(
        \pk_indw_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9554 ), .A(
        \SADR/ADDIDX/add_w_x_z/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9556 ), .A(\SADR/pgaddxz[14] ), .B(
        \pk_indw_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9558 ), .A(\SADR/pgaddxz[15] ), .B(
        \pk_indw_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add2/n9549 ), .A(
        \SADR/ADDIDX/add_w_x_z/add2/n9548 ), .B(
        \SADR/ADDIDX/add_w_x_z/add2/n9529 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/c_last ), .A(\SADR/ADDIDX/add_w_x_z/add3/n9495 
        ), .B(\SADR/ADDIDX/add_w_x_z/add3/n9496 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9497 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/gp_out[3] ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9498 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9495 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9499 ), .D(
        \SADR/ADDIDX/add_w_x_z/add3/n9500 ), .E(
        \SADR/ADDIDX/add_w_x_z/add3/n9501 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9511 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9510 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9512 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add3/n9513 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9498 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9514 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9514 ), .A(\SADR/pgaddxz[18] ), .B(
        \pk_indw_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9516 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9495 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9509 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9512 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9498 ), .A(\SADR/pgaddxz[18] ), .B(
        \pk_indw_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9497 ), .A(\SADR/pgaddxz[22] ), .B(
        \pk_indw_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9519 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9520 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9524 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add3/U26  ( .Z(\SADR/pgaddwxz[18] ), .A(
        \SADR/ADDIDX/add_w_x_z/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9513 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_z/gg_out[3] ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9501 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9502 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9503 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9507 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9508 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9509 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9510 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9518 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9522 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9498 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9500 ), .D(
        \SADR/ADDIDX/add_w_x_z/add3/n9523 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9495 ), .A(\SADR/pgaddxz[22] ), .B(
        \pk_indw_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9496 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9518 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9525 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9506 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add3/U20  ( .Z(\SADR/pgaddwxz[19] ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9508 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9511 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9520 ), .A(\SADR/pgaddxz[20] ), .B(
        \pk_indw_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9515 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9523 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9499 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9526 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9504 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9503 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9501 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9502 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9515 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9516 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9497 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add3/U17  ( .Z(\SADR/pgaddwxz[22] ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9517 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9496 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9500 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9520 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9509 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9512 ), .A(\SADR/pgaddxz[19] ), .B(
        \pk_indw_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9506 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9526 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9510 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9521 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9501 ), .A(\SADR/pgaddxz[23] ), .B(
        \pk_indw_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9508 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9498 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9522 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9514 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9505 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9506 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9499 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add3/U19  ( .Z(\SADR/pgaddwxz[20] ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9519 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9507 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add3/n9523 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9514 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9500 ), .C(
        \SADR/ADDIDX/add_w_x_z/add3/n9520 ), .D(
        \SADR/ADDIDX/add_w_x_z/add3/n9521 ), .E(
        \SADR/ADDIDX/add_w_x_z/add3/n9524 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9525 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9499 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add3/U16  ( .Z(\SADR/pgaddwxz[23] ), .A(
        \SADR/ADDIDX/add_w_x_z/c_last ), .B(\SADR/ADDIDX/add_w_x_z/add3/n9504 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_z/add3/U18  ( .Z(\SADR/pgaddwxz[21] ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9518 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9505 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9499 ), .A(\SADR/pgaddxz[21] ), .B(
        \pk_indw_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_z/add3/n9503 ), .A(\SADR/pgaddxz[23] ), .B(
        \pk_indw_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9521 ), .A(\SADR/pgaddxz[19] ), .B(
        \pk_indw_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9522 ), .A(
        \SADR/ADDIDX/add_w_x_z/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9524 ), .A(\SADR/pgaddxz[20] ), .B(
        \pk_indw_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9526 ), .A(\SADR/pgaddxz[21] ), .B(
        \pk_indw_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_z/add3/n9517 ), .A(
        \SADR/ADDIDX/add_w_x_z/add3/n9516 ), .B(
        \SADR/ADDIDX/add_w_x_z/add3/n9497 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9462 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9463 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9464 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9465 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9462 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9466 ), .D(
        \SADR/ADDIDX/add_w_y_z/add0/n9467 ), .E(
        \SADR/ADDIDX/add_w_y_z/add0/n9468 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9478 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9477 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9479 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add0/n9480 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9465 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9481 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9481 ), .A(\SADR/pgaddwy[0] ), .B(
        \pk_indz_h[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9483 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9462 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9476 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9479 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9465 ), .A(\SADR/pgaddwy[0] ), .B(
        \pk_indz_h[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9464 ), .A(\SADR/pgaddwy[4] ), .B(
        \pk_indz_h[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9486 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9487 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9491 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add0/U26  ( .Z(\SADR/pgaddwyz[0] ), .A(
        1'b0), .B(\SADR/ADDIDX/add_w_y_z/add0/n9480 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_y_z/gg_out[0] ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9468 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9469 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9470 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9474 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9475 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9476 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9477 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9485 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9489 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9465 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9467 ), .D(
        \SADR/ADDIDX/add_w_y_z/add0/n9490 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9462 ), .A(\SADR/pgaddwy[4] ), .B(
        \pk_indz_h[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9463 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9485 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9492 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9473 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add0/U20  ( .Z(\SADR/pgaddwyz[1] ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9475 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9478 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9487 ), .A(\SADR/pgaddwy[2] ), .B(
        \pk_indz_h[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9482 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9490 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9466 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9493 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9471 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9470 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9468 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9469 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9482 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9483 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9464 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add0/U17  ( .Z(\SADR/pgaddwyz[4] ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9484 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9463 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9467 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9487 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9476 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9479 ), .A(\SADR/pgaddwy[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9473 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9493 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9477 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9488 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9468 ), .A(\SADR/pgaddwy[5] ), .B(
        \pk_indz_h[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9475 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9465 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9489 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9481 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9472 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9473 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9466 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add0/U19  ( .Z(\SADR/pgaddwyz[2] ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9486 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9474 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add0/n9490 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9481 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9467 ), .C(
        \SADR/ADDIDX/add_w_y_z/add0/n9487 ), .D(
        \SADR/ADDIDX/add_w_y_z/add0/n9488 ), .E(
        \SADR/ADDIDX/add_w_y_z/add0/n9491 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9492 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9466 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add0/U16  ( .Z(\SADR/pgaddwyz[5] ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9471 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add0/U18  ( .Z(\SADR/pgaddwyz[3] ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9485 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9472 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9466 ), .A(\SADR/pgaddwy[3] ), .B(
        \pk_indz_h[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add0/n9470 ), .A(\SADR/pgaddwy[5] ), .B(
        \pk_indz_h[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9488 ), .A(\SADR/pgaddwy[1] ), .B(
        \pk_indz_h[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9489 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9491 ), .A(\SADR/pgaddwy[2] ), .B(
        \pk_indz_h[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9493 ), .A(\SADR/pgaddwy[3] ), .B(
        \pk_indz_h[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add0/n9484 ), .A(
        \SADR/ADDIDX/add_w_y_z/add0/n9483 ), .B(
        \SADR/ADDIDX/add_w_y_z/add0/n9464 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9430 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9431 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9432 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/gp_out[1] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9433 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9430 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9434 ), .D(
        \SADR/ADDIDX/add_w_y_z/add1/n9435 ), .E(
        \SADR/ADDIDX/add_w_y_z/add1/n9436 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9446 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9445 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9447 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add1/n9448 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9433 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9449 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9449 ), .A(\SADR/pgaddwy[6] ), .B(
        \pk_indz_h[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9451 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9430 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9444 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9447 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9433 ), .A(\SADR/pgaddwy[6] ), .B(
        \pk_indz_h[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9432 ), .A(\SADR/pgaddwy[10] ), .B(
        \pk_indz_h[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9454 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9455 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9459 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add1/U26  ( .Z(\SADR/pgaddwyz[6] ), .A(
        \SADR/ADDIDX/add_w_y_z/gg_out[0] ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9448 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_y_z/gg_out[1] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9436 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9437 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9438 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9442 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9443 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9444 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9445 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9453 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9457 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9433 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9435 ), .D(
        \SADR/ADDIDX/add_w_y_z/add1/n9458 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9430 ), .A(\SADR/pgaddwy[10] ), .B(
        \pk_indz_h[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9431 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9453 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9460 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9441 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add1/U20  ( .Z(\SADR/pgaddwyz[7] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9443 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9446 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9455 ), .A(\SADR/pgaddwy[8] ), .B(
        \pk_indz_h[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9450 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9458 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9434 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9461 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9439 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9438 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9436 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9437 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9450 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9451 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9432 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add1/U17  ( .Z(\SADR/pgaddwyz[10] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9452 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9431 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9435 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9455 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9444 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9447 ), .A(\SADR/pgaddwy[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9441 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9461 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9445 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9456 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9436 ), .A(\SADR/pgaddwy[11] ), .B(
        \pk_indz_h[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9443 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9433 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9457 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9449 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9440 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9441 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9434 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add1/U19  ( .Z(\SADR/pgaddwyz[8] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9454 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9442 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add1/n9458 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9449 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9435 ), .C(
        \SADR/ADDIDX/add_w_y_z/add1/n9455 ), .D(
        \SADR/ADDIDX/add_w_y_z/add1/n9456 ), .E(
        \SADR/ADDIDX/add_w_y_z/add1/n9459 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9460 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9434 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add1/U16  ( .Z(\SADR/pgaddwyz[11] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9439 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add1/U18  ( .Z(\SADR/pgaddwyz[9] ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9453 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9440 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9434 ), .A(\SADR/pgaddwy[9] ), .B(
        \pk_indz_h[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add1/n9438 ), .A(\SADR/pgaddwy[11] ), .B(
        \pk_indz_h[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9456 ), .A(\SADR/pgaddwy[7] ), .B(
        \pk_indz_h[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9457 ), .A(
        \SADR/ADDIDX/add_w_y_z/gg_out[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9459 ), .A(\SADR/pgaddwy[8] ), .B(
        \pk_indz_h[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9461 ), .A(\SADR/pgaddwy[9] ), .B(
        \pk_indz_h[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add1/n9452 ), .A(
        \SADR/ADDIDX/add_w_y_z/add1/n9451 ), .B(
        \SADR/ADDIDX/add_w_y_z/add1/n9432 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9398 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9399 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9400 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/gp_out[2] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9401 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9398 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9402 ), .D(
        \SADR/ADDIDX/add_w_y_z/add2/n9403 ), .E(
        \SADR/ADDIDX/add_w_y_z/add2/n9404 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9414 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9413 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9415 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add2/n9416 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9401 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9417 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9417 ), .A(\SADR/pgaddwy[12] ), .B(
        \pk_indz_h[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9419 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9398 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9412 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9415 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9401 ), .A(\SADR/pgaddwy[12] ), .B(
        \pk_indz_h[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9400 ), .A(\SADR/pgaddwy[16] ), .B(
        \pk_indz_h[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9422 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9423 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9427 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add2/U26  ( .Z(\SADR/pgaddwyz[12] ), .A(
        \SADR/ADDIDX/add_w_y_z/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9416 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_y_z/gg_out[2] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9404 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9405 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9406 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9410 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9411 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9412 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9413 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9421 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9425 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9401 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9403 ), .D(
        \SADR/ADDIDX/add_w_y_z/add2/n9426 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9398 ), .A(\SADR/pgaddwy[16] ), .B(
        \pk_indz_h[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9399 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9421 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9428 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9409 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add2/U20  ( .Z(\SADR/pgaddwyz[13] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9411 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9414 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9423 ), .A(\SADR/pgaddwy[14] ), .B(
        \pk_indz_h[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9418 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9426 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9402 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9429 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9407 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9406 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9404 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9405 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9418 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9419 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9400 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add2/U17  ( .Z(\SADR/pgaddwyz[16] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9420 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9399 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9403 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9423 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9412 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9415 ), .A(\SADR/pgaddwy[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9409 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9429 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9413 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9424 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9404 ), .A(\SADR/pgaddwy[17] ), .B(
        \pk_indz_h[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9411 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9401 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9425 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9417 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9408 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9409 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9402 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add2/U19  ( .Z(\SADR/pgaddwyz[14] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9422 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9410 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add2/n9426 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9417 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9403 ), .C(
        \SADR/ADDIDX/add_w_y_z/add2/n9423 ), .D(
        \SADR/ADDIDX/add_w_y_z/add2/n9424 ), .E(
        \SADR/ADDIDX/add_w_y_z/add2/n9427 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9428 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9402 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add2/U16  ( .Z(\SADR/pgaddwyz[17] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9407 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add2/U18  ( .Z(\SADR/pgaddwyz[15] ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9421 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9408 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9402 ), .A(\SADR/pgaddwy[15] ), .B(
        \pk_indz_h[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add2/n9406 ), .A(\SADR/pgaddwy[17] ), .B(
        \pk_indz_h[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9424 ), .A(\SADR/pgaddwy[13] ), .B(
        \pk_indz_h[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9425 ), .A(
        \SADR/ADDIDX/add_w_y_z/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9427 ), .A(\SADR/pgaddwy[14] ), .B(
        \pk_indz_h[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9429 ), .A(\SADR/pgaddwy[15] ), .B(
        \pk_indz_h[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add2/n9420 ), .A(
        \SADR/ADDIDX/add_w_y_z/add2/n9419 ), .B(
        \SADR/ADDIDX/add_w_y_z/add2/n9400 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/c_last ), .A(\SADR/ADDIDX/add_w_y_z/add3/n9366 
        ), .B(\SADR/ADDIDX/add_w_y_z/add3/n9367 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9368 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_y_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/gp_out[3] ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9369 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9366 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9370 ), .D(
        \SADR/ADDIDX/add_w_y_z/add3/n9371 ), .E(
        \SADR/ADDIDX/add_w_y_z/add3/n9372 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9382 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9381 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9383 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_y_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add3/n9384 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9369 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9385 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9385 ), .A(\SADR/pgaddwy[18] ), .B(
        \pk_indz_h[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9387 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9366 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9380 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9383 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9369 ), .A(\SADR/pgaddwy[18] ), .B(
        \pk_indz_h[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9368 ), .A(\SADR/pgaddwy[22] ), .B(
        \pk_indz_h[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9390 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9391 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9395 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add3/U26  ( .Z(\SADR/pgaddwyz[18] ), .A(
        \SADR/ADDIDX/add_w_y_z/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9384 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_y_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_y_z/gg_out[3] ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9372 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9373 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9374 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9378 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9379 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9380 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9381 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_y_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9389 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9393 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9369 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9371 ), .D(
        \SADR/ADDIDX/add_w_y_z/add3/n9394 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9366 ), .A(\SADR/pgaddwy[22] ), .B(
        \pk_indz_h[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_y_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9367 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9389 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9396 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9377 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add3/U20  ( .Z(\SADR/pgaddwyz[19] ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9379 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9382 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9391 ), .A(\SADR/pgaddwy[20] ), .B(
        \pk_indz_h[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9386 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9394 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9370 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9397 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9375 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9374 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9372 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_y_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9373 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9386 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9387 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9368 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add3/U17  ( .Z(\SADR/pgaddwyz[22] ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9388 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9367 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_y_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9371 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9391 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9380 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9383 ), .A(\SADR/pgaddwy[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9377 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9397 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9381 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9392 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9372 ), .A(\SADR/pgaddwy[23] ), .B(
        \pk_indz_h[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_y_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9379 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9369 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9393 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9385 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9376 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9377 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9370 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add3/U19  ( .Z(\SADR/pgaddwyz[20] ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9390 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9378 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_y_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add3/n9394 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9385 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9371 ), .C(
        \SADR/ADDIDX/add_w_y_z/add3/n9391 ), .D(
        \SADR/ADDIDX/add_w_y_z/add3/n9392 ), .E(
        \SADR/ADDIDX/add_w_y_z/add3/n9395 ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9396 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9370 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add3/U16  ( .Z(\SADR/pgaddwyz[23] ), .A(
        \SADR/ADDIDX/add_w_y_z/c_last ), .B(\SADR/ADDIDX/add_w_y_z/add3/n9375 
        ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_y_z/add3/U18  ( .Z(\SADR/pgaddwyz[21] ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9389 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9376 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_y_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9370 ), .A(\SADR/pgaddwy[21] ), .B(
        \pk_indz_h[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_y_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_y_z/add3/n9374 ), .A(\SADR/pgaddwy[23] ), .B(
        \pk_indz_h[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9392 ), .A(\SADR/pgaddwy[19] ), .B(
        \pk_indz_h[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_y_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9393 ), .A(
        \SADR/ADDIDX/add_w_y_z/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9395 ), .A(\SADR/pgaddwy[20] ), .B(
        \pk_indz_h[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9397 ), .A(\SADR/pgaddwy[21] ), .B(
        \pk_indz_h[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_y_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_y_z/add3/n9388 ), .A(
        \SADR/ADDIDX/add_w_y_z/add3/n9387 ), .B(
        \SADR/ADDIDX/add_w_y_z/add3/n9368 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add0/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9333 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9334 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9335 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y_z/add0/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/gp_out ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9336 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9333 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9337 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9338 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9339 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9349 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9348 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9350 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y_z/add0/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9351 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9336 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9352 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9352 ), .A(\SADR/pgaddwz[0] ), .B(
        \SADR/pgaddxy[0] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add0/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9354 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9333 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add0/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9347 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9350 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9336 ), .A(\SADR/pgaddwz[0] ), .B(
        \SADR/pgaddxy[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9335 ), .A(\SADR/pgaddwz[4] ), .B(
        \SADR/pgaddxy[4] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add0/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9357 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9358 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9362 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U26  ( .Z(\SADR/pgaddwxyz[0] ), 
        .A(1'b0), .B(\SADR/ADDIDX/add_w_x_y_z/add0/n9351 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[0] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9339 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9340 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9341 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add0/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9345 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9346 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9347 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9348 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y_z/add0/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9356 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9360 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9336 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9338 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9361 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9333 ), .A(\SADR/pgaddwz[4] ), .B(
        \SADR/pgaddxy[4] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add0/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9334 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9356 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9363 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9344 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U20  ( .Z(\SADR/pgaddwxyz[1] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add0/n9346 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9349 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9358 ), .A(\SADR/pgaddwz[2] ), .B(
        \SADR/pgaddxy[2] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add0/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9353 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9361 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9337 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9364 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9342 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9341 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9339 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y_z/add0/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9340 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9353 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9354 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9335 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U17  ( .Z(\SADR/pgaddwxyz[4] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add0/n9355 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9334 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add0/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9338 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9358 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9347 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9350 ), .A(\SADR/pgaddwz[1] ), .B(
        \SADR/pgaddxy[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add0/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9344 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9364 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add0/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9348 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9359 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9339 ), .A(\SADR/pgaddwz[5] ), .B(
        \SADR/pgaddxy[5] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add0/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9346 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9336 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9360 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9352 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9343 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9344 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9337 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U19  ( .Z(\SADR/pgaddwxyz[2] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add0/n9357 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9345 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y_z/add0/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9361 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9352 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9338 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9358 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9359 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9362 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add0/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9363 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9337 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U16  ( .Z(\SADR/pgaddwxyz[5] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add0/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9342 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add0/U18  ( .Z(\SADR/pgaddwxyz[3] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add0/n9356 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9343 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9337 ), .A(\SADR/pgaddwz[3] ), .B(
        \SADR/pgaddxy[3] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9341 ), .A(\SADR/pgaddwz[5] ), .B(
        \SADR/pgaddxy[5] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9359 ), .A(\SADR/pgaddwz[1] ), .B(
        \SADR/pgaddxy[1] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add0/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9360 ), .A(1'b0) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9362 ), .A(\SADR/pgaddwz[2] ), .B(
        \SADR/pgaddxy[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9364 ), .A(\SADR/pgaddwz[3] ), .B(
        \SADR/pgaddxy[3] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add0/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9355 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9354 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add0/n9335 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add1/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9301 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9302 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9303 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y_z/add1/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/gp_out[1] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9304 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9301 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9305 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9306 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9307 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9317 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9316 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9318 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y_z/add1/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9319 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9304 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9320 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9320 ), .A(\SADR/pgaddwz[6] ), .B(
        \SADR/pgaddxy[6] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add1/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9322 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9301 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add1/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9315 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9318 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9304 ), .A(\SADR/pgaddwz[6] ), .B(
        \SADR/pgaddxy[6] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9303 ), .A(\SADR/pgaddwz[10] ), .B(
        \SADR/pgaddxy[10] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add1/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9325 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9326 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9330 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U26  ( .Z(\SADR/pgaddwxyz[6] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/gg_out[0] ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9319 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[1] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9307 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9308 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9309 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add1/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9313 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9314 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9315 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9316 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y_z/add1/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9324 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9328 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9304 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9306 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9329 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9301 ), .A(\SADR/pgaddwz[10] ), .B(
        \SADR/pgaddxy[10] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add1/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9302 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9324 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9331 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9312 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U20  ( .Z(\SADR/pgaddwxyz[7] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add1/n9314 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9317 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9326 ), .A(\SADR/pgaddwz[8] ), .B(
        \SADR/pgaddxy[8] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add1/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9321 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9329 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9305 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9332 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9310 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9309 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9307 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y_z/add1/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9308 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9321 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9322 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9303 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U17  ( .Z(\SADR/pgaddwxyz[10] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add1/n9323 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9302 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add1/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9306 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9326 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9315 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9318 ), .A(\SADR/pgaddwz[7] ), .B(
        \SADR/pgaddxy[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add1/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9312 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9332 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add1/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9316 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9327 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9307 ), .A(\SADR/pgaddwz[11] ), .B(
        \SADR/pgaddxy[11] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add1/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9314 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9304 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9328 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9320 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9311 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9312 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9305 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U19  ( .Z(\SADR/pgaddwxyz[8] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add1/n9325 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9313 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y_z/add1/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9329 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9320 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9306 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9326 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9327 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9330 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add1/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9331 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9305 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U16  ( .Z(\SADR/pgaddwxyz[11] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add1/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9310 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add1/U18  ( .Z(\SADR/pgaddwxyz[9] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add1/n9324 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9311 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9305 ), .A(\SADR/pgaddwz[9] ), .B(
        \SADR/pgaddxy[9] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9309 ), .A(\SADR/pgaddwz[11] ), .B(
        \SADR/pgaddxy[11] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9327 ), .A(\SADR/pgaddwz[7] ), .B(
        \SADR/pgaddxy[7] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add1/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9328 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[0] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9330 ), .A(\SADR/pgaddwz[8] ), .B(
        \SADR/pgaddxy[8] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9332 ), .A(\SADR/pgaddwz[9] ), .B(
        \SADR/pgaddxy[9] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add1/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9323 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9322 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add1/n9303 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add2/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9269 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9270 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9271 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y_z/add2/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/gp_out[2] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9272 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9269 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9273 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9274 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9275 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9285 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9284 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9286 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y_z/add2/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9287 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9272 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9288 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9288 ), .A(\SADR/pgaddwz[12] ), .B(
        \SADR/pgaddxy[12] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add2/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9290 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9269 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add2/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9283 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9286 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9272 ), .A(\SADR/pgaddwz[12] ), .B(
        \SADR/pgaddxy[12] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9271 ), .A(\SADR/pgaddwz[16] ), .B(
        \SADR/pgaddxy[16] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add2/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9293 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9294 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9298 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U26  ( .Z(\SADR/pgaddwxyz[12] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/cin_stg[1] ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9287 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[2] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9275 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9276 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9277 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add2/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9281 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9282 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9283 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9284 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y_z/add2/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9292 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9296 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9272 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9274 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9297 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9269 ), .A(\SADR/pgaddwz[16] ), .B(
        \SADR/pgaddxy[16] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add2/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9270 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9292 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9299 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9280 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U20  ( .Z(\SADR/pgaddwxyz[13] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add2/n9282 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9285 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9294 ), .A(\SADR/pgaddwz[14] ), .B(
        \SADR/pgaddxy[14] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add2/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9289 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9297 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9273 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9300 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9278 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9277 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9275 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y_z/add2/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9276 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9289 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9290 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9271 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U17  ( .Z(\SADR/pgaddwxyz[16] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add2/n9291 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9270 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add2/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9274 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9294 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9283 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9286 ), .A(\SADR/pgaddwz[13] ), .B(
        \SADR/pgaddxy[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add2/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9280 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9300 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add2/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9284 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9295 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9275 ), .A(\SADR/pgaddwz[17] ), .B(
        \SADR/pgaddxy[17] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add2/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9282 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9272 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9296 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9288 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9279 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9280 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9273 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U19  ( .Z(\SADR/pgaddwxyz[14] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add2/n9293 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9281 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y_z/add2/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9297 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9288 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9274 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9294 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9295 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9298 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add2/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9299 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9273 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U16  ( .Z(\SADR/pgaddwxyz[17] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add2/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9278 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add2/U18  ( .Z(\SADR/pgaddwxyz[15] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add2/n9292 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9279 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9273 ), .A(\SADR/pgaddwz[15] ), .B(
        \SADR/pgaddxy[15] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9277 ), .A(\SADR/pgaddwz[17] ), .B(
        \SADR/pgaddxy[17] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9295 ), .A(\SADR/pgaddwz[13] ), .B(
        \SADR/pgaddxy[13] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add2/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9296 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[1] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9298 ), .A(\SADR/pgaddwz[14] ), .B(
        \SADR/pgaddxy[14] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9300 ), .A(\SADR/pgaddwz[15] ), .B(
        \SADR/pgaddxy[15] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add2/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9291 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9290 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add2/n9271 ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add3/U7  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/c_last ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9237 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9238 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9239 ) );
    snl_nor05x1 \SADR/ADDIDX/add_w_x_y_z/add3/U8  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/gp_out[3] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9240 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9237 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9241 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9242 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9243 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U13  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9253 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9252 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9254 ) );
    snl_and12x1 \SADR/ADDIDX/add_w_x_y_z/add3/U14  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9255 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9240 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9256 ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U21  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9256 ), .A(\SADR/pgaddwz[18] ), .B(
        \SADR/pgaddxy[18] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add3/U28  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9258 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9237 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add3/U33  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9251 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9254 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U34  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9240 ), .A(\SADR/pgaddwz[18] ), .B(
        \SADR/pgaddxy[18] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U41  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9239 ), .A(\SADR/pgaddwz[22] ), .B(
        \SADR/pgaddxy[22] ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add3/U46  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9261 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9262 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9266 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U26  ( .Z(\SADR/pgaddwxyz[18] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/cin_stg[2] ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9255 ) );
    snl_ao01b2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U9  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/gg_out[3] ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9243 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9244 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9245 ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add3/U12  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9249 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9250 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9251 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9252 ) );
    snl_oai013x0 \SADR/ADDIDX/add_w_x_y_z/add3/U35  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9260 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9264 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9240 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9242 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9265 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U27  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9237 ), .A(\SADR/pgaddwz[22] ), .B(
        \SADR/pgaddxy[22] ) );
    snl_aoi012x1 \SADR/ADDIDX/add_w_x_y_z/add3/U40  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9238 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9260 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9267 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9248 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U20  ( .Z(\SADR/pgaddwxyz[19] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add3/n9250 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9253 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U29  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9262 ), .A(\SADR/pgaddwz[20] ), .B(
        \SADR/pgaddxy[20] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add3/U47  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9257 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9265 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9241 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9268 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U10  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9246 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9245 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9243 ) );
    snl_aoi0b12x0 \SADR/ADDIDX/add_w_x_y_z/add3/U15  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9244 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9257 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9258 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9239 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U17  ( .Z(\SADR/pgaddwxyz[22] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add3/n9259 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9238 ) );
    snl_nand12x1 \SADR/ADDIDX/add_w_x_y_z/add3/U22  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9242 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9262 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9251 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U32  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9254 ), .A(\SADR/pgaddwz[19] ), .B(
        \SADR/pgaddxy[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add3/U39  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9248 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9268 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add3/U30  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9252 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9263 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U42  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9243 ), .A(\SADR/pgaddwz[23] ), .B(
        \SADR/pgaddxy[23] ) );
    snl_oai012x1 \SADR/ADDIDX/add_w_x_y_z/add3/U45  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9250 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9240 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9264 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9256 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U11  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9247 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9248 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9241 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U19  ( .Z(\SADR/pgaddwxyz[20] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add3/n9261 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9249 ) );
    snl_oa122x1 \SADR/ADDIDX/add_w_x_y_z/add3/U25  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9265 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9256 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9242 ), .C(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9262 ), .D(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9263 ), .E(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9266 ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add3/U37  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9267 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9241 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U16  ( .Z(\SADR/pgaddwxyz[23] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/c_last ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9246 ) );
    snl_xor2x0 \SADR/ADDIDX/add_w_x_y_z/add3/U18  ( .Z(\SADR/pgaddwxyz[21] ), 
        .A(\SADR/ADDIDX/add_w_x_y_z/add3/n9260 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9247 ) );
    snl_nor02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U36  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9241 ), .A(\SADR/pgaddwz[21] ), .B(
        \SADR/pgaddxy[21] ) );
    snl_and02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U43  ( .Z(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9245 ), .A(\SADR/pgaddwz[23] ), .B(
        \SADR/pgaddxy[23] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U23  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9263 ), .A(\SADR/pgaddwz[19] ), .B(
        \SADR/pgaddxy[19] ) );
    snl_invx05 \SADR/ADDIDX/add_w_x_y_z/add3/U24  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9264 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/cin_stg[2] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U31  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9266 ), .A(\SADR/pgaddwz[20] ), .B(
        \SADR/pgaddxy[20] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U38  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9268 ), .A(\SADR/pgaddwz[21] ), .B(
        \SADR/pgaddxy[21] ) );
    snl_nand02x1 \SADR/ADDIDX/add_w_x_y_z/add3/U44  ( .ZN(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9259 ), .A(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9258 ), .B(
        \SADR/ADDIDX/add_w_x_y_z/add3/n9239 ) );
    snl_ao012x1 \REGF/pbmemff41/phdec12_2/dec4_1/U7  ( .Z(
        \REGF/pbmemff41/RO_TRCOT[0] ), .A(\pk_stdat[0] ), .B(1'b0), .C(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7075 ) );
    snl_or04x1 \REGF/pbmemff41/phdec12_2/dec4_1/U8  ( .Z(
        \REGF/pbmemff41/phdec12_2/gg_out[0] ), .A(\pk_stdat[0] ), .B(
        \pk_stdat[3] ), .C(\pk_stdat[1] ), .D(\pk_stdat[2] ) );
    snl_nand02x1 \REGF/pbmemff41/phdec12_2/dec4_1/U13  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7079 ), .A(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7075 ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7078 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_2/dec4_1/U14  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7077 ), .A(\pk_stdat[3] ) );
    snl_oai022x1 \REGF/pbmemff41/phdec12_2/dec4_1/U9  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[3] ), .A(1'b0), .B(
        \REGF/pbmemff41/phdec12_2/gg_out[0] ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7076 ), .D(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7077 ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_2/dec4_1/U12  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7075 ), .A(1'b0), .B(\pk_stdat[0] )
         );
    snl_oai012x1 \REGF/pbmemff41/phdec12_2/dec4_1/U10  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[1] ), .A(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7075 ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7078 ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7079 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_2/dec4_1/U15  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7078 ), .A(\pk_stdat[1] ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_2/dec4_1/U11  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7076 ), .A(\pk_stdat[2] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7079 ) );
    snl_xnor2x0 \REGF/pbmemff41/phdec12_2/dec4_1/U16  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[2] ), .A(\pk_stdat[2] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_1/n7079 ) );
    snl_ao012x1 \REGF/pbmemff41/phdec12_2/dec4_3/U7  ( .Z(
        \REGF/pbmemff41/RO_TRCOT[8] ), .A(\pk_stdat[8] ), .B(
        \REGF/pbmemff41/phdec12_2/gcarry[1] ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7070 ) );
    snl_or04x1 \REGF/pbmemff41/phdec12_2/dec4_3/U8  ( .Z(
        \REGF/pbmemff41/phdec12_2/dec4_3/gg_out ), .A(\pk_stdat[8] ), .B(
        \pk_stdat[11] ), .C(\pk_stdat[9] ), .D(\pk_stdat[10] ) );
    snl_nand02x1 \REGF/pbmemff41/phdec12_2/dec4_3/U13  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7074 ), .A(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7070 ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7073 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_2/dec4_3/U14  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7072 ), .A(\pk_stdat[11] ) );
    snl_oai022x1 \REGF/pbmemff41/phdec12_2/dec4_3/U9  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[11] ), .A(
        \REGF/pbmemff41/phdec12_2/gcarry[1] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_3/gg_out ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7071 ), .D(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7072 ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_2/dec4_3/U12  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7070 ), .A(
        \REGF/pbmemff41/phdec12_2/gcarry[1] ), .B(\pk_stdat[8] ) );
    snl_oai012x1 \REGF/pbmemff41/phdec12_2/dec4_3/U10  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[9] ), .A(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7070 ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7073 ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7074 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_2/dec4_3/U15  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7073 ), .A(\pk_stdat[9] ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_2/dec4_3/U11  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7071 ), .A(\pk_stdat[10] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7074 ) );
    snl_xnor2x0 \REGF/pbmemff41/phdec12_2/dec4_3/U16  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[10] ), .A(\pk_stdat[10] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_3/n7074 ) );
    snl_ao012x1 \REGF/pbmemff41/phdec12_2/dec4_2/U7  ( .Z(
        \REGF/pbmemff41/RO_TRCOT[4] ), .A(\pk_stdat[4] ), .B(
        \REGF/pbmemff41/phdec12_2/gg_out[0] ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7065 ) );
    snl_or04x1 \REGF/pbmemff41/phdec12_2/dec4_2/U8  ( .Z(
        \REGF/pbmemff41/phdec12_2/gg_out[1] ), .A(\pk_stdat[4] ), .B(
        \pk_stdat[7] ), .C(\pk_stdat[5] ), .D(\pk_stdat[6] ) );
    snl_nand02x1 \REGF/pbmemff41/phdec12_2/dec4_2/U13  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7069 ), .A(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7065 ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7068 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_2/dec4_2/U14  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7067 ), .A(\pk_stdat[7] ) );
    snl_oai022x1 \REGF/pbmemff41/phdec12_2/dec4_2/U9  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[7] ), .A(\REGF/pbmemff41/phdec12_2/gg_out[0] 
        ), .B(\REGF/pbmemff41/phdec12_2/gg_out[1] ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7066 ), .D(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7067 ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_2/dec4_2/U12  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7065 ), .A(
        \REGF/pbmemff41/phdec12_2/gg_out[0] ), .B(\pk_stdat[4] ) );
    snl_oai012x1 \REGF/pbmemff41/phdec12_2/dec4_2/U10  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[5] ), .A(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7065 ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7068 ), .C(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7069 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_2/dec4_2/U15  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7068 ), .A(\pk_stdat[5] ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_2/dec4_2/U11  ( .ZN(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7066 ), .A(\pk_stdat[6] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7069 ) );
    snl_xnor2x0 \REGF/pbmemff41/phdec12_2/dec4_2/U16  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[6] ), .A(\pk_stdat[6] ), .B(
        \REGF/pbmemff41/phdec12_2/dec4_2/n7069 ) );
    snl_ao012x1 \REGF/pbmemff41/phdec12_1/dec4_1/U7  ( .Z(
        \REGF/pbmemff41/RO_TRCOT[12] ), .A(\pk_stdat[12] ), .B(1'b0), .C(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7058 ) );
    snl_or04x1 \REGF/pbmemff41/phdec12_1/dec4_1/U8  ( .Z(
        \REGF/pbmemff41/phdec12_1/gg_out[0] ), .A(\pk_stdat[12] ), .B(
        \pk_stdat[15] ), .C(\pk_stdat[13] ), .D(\pk_stdat[14] ) );
    snl_nand02x1 \REGF/pbmemff41/phdec12_1/dec4_1/U13  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7062 ), .A(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7058 ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7061 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_1/dec4_1/U14  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7060 ), .A(\pk_stdat[15] ) );
    snl_oai022x1 \REGF/pbmemff41/phdec12_1/dec4_1/U9  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[15] ), .A(1'b0), .B(
        \REGF/pbmemff41/phdec12_1/gg_out[0] ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7059 ), .D(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7060 ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_1/dec4_1/U12  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7058 ), .A(1'b0), .B(\pk_stdat[12] )
         );
    snl_oai012x1 \REGF/pbmemff41/phdec12_1/dec4_1/U10  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[13] ), .A(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7058 ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7061 ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7062 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_1/dec4_1/U15  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7061 ), .A(\pk_stdat[13] ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_1/dec4_1/U11  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7059 ), .A(\pk_stdat[14] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7062 ) );
    snl_xnor2x0 \REGF/pbmemff41/phdec12_1/dec4_1/U16  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[14] ), .A(\pk_stdat[14] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_1/n7062 ) );
    snl_ao012x1 \REGF/pbmemff41/phdec12_1/dec4_3/U7  ( .Z(
        \REGF/pbmemff41/RO_TRCOT[20] ), .A(\pk_stdat[20] ), .B(
        \REGF/pbmemff41/phdec12_1/gcarry[1] ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7053 ) );
    snl_or04x1 \REGF/pbmemff41/phdec12_1/dec4_3/U8  ( .Z(
        \REGF/pbmemff41/phdec12_1/dec4_3/gg_out ), .A(\pk_stdat[20] ), .B(
        \REGF/RO_TRCO[27] ), .C(\REGF/RO_TRCO[25] ), .D(\REGF/RO_TRCO[26] ) );
    snl_nand02x1 \REGF/pbmemff41/phdec12_1/dec4_3/U13  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7057 ), .A(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7053 ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7056 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_1/dec4_3/U14  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7055 ), .A(\REGF/RO_TRCO[27] ) );
    snl_oai022x1 \REGF/pbmemff41/phdec12_1/dec4_3/U9  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[23] ), .A(
        \REGF/pbmemff41/phdec12_1/gcarry[1] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_3/gg_out ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7054 ), .D(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7055 ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_1/dec4_3/U12  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7053 ), .A(
        \REGF/pbmemff41/phdec12_1/gcarry[1] ), .B(\pk_stdat[20] ) );
    snl_oai012x1 \REGF/pbmemff41/phdec12_1/dec4_3/U10  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[21] ), .A(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7053 ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7056 ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7057 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_1/dec4_3/U15  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7056 ), .A(\REGF/RO_TRCO[25] ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_1/dec4_3/U11  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7054 ), .A(\REGF/RO_TRCO[26] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7057 ) );
    snl_xnor2x0 \REGF/pbmemff41/phdec12_1/dec4_3/U16  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[22] ), .A(\REGF/RO_TRCO[26] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_3/n7057 ) );
    snl_ao012x1 \REGF/pbmemff41/phdec12_1/dec4_2/U7  ( .Z(
        \REGF/pbmemff41/RO_TRCOT[16] ), .A(\pk_stdat[16] ), .B(
        \REGF/pbmemff41/phdec12_1/gg_out[0] ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7048 ) );
    snl_or04x1 \REGF/pbmemff41/phdec12_1/dec4_2/U8  ( .Z(
        \REGF/pbmemff41/phdec12_1/gg_out[1] ), .A(\pk_stdat[16] ), .B(
        \pk_stdat[19] ), .C(\pk_stdat[17] ), .D(\pk_stdat[18] ) );
    snl_nand02x1 \REGF/pbmemff41/phdec12_1/dec4_2/U13  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7052 ), .A(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7048 ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7051 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_1/dec4_2/U14  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7050 ), .A(\pk_stdat[19] ) );
    snl_oai022x1 \REGF/pbmemff41/phdec12_1/dec4_2/U9  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[19] ), .A(
        \REGF/pbmemff41/phdec12_1/gg_out[0] ), .B(
        \REGF/pbmemff41/phdec12_1/gg_out[1] ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7049 ), .D(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7050 ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_1/dec4_2/U12  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7048 ), .A(
        \REGF/pbmemff41/phdec12_1/gg_out[0] ), .B(\pk_stdat[16] ) );
    snl_oai012x1 \REGF/pbmemff41/phdec12_1/dec4_2/U10  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[17] ), .A(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7048 ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7051 ), .C(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7052 ) );
    snl_invx05 \REGF/pbmemff41/phdec12_1/dec4_2/U15  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7051 ), .A(\pk_stdat[17] ) );
    snl_nor02x1 \REGF/pbmemff41/phdec12_1/dec4_2/U11  ( .ZN(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7049 ), .A(\pk_stdat[18] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7052 ) );
    snl_xnor2x0 \REGF/pbmemff41/phdec12_1/dec4_2/U16  ( .ZN(
        \REGF/pbmemff41/RO_TRCOT[18] ), .A(\pk_stdat[18] ), .B(
        \REGF/pbmemff41/phdec12_1/dec4_2/n7052 ) );
    snl_aoi112x0 \MAIN/ENGIN/STEP_A/deocgen_1/U12  ( .ZN(
        \MAIN/ENGIN/a_deocenh ), .A(\MAIN/ENGIN/STEP_A/cst[0] ), .B(
        \MAIN/ENGIN/STEP_A/deocgen_1/n3543 ), .C(\MAIN/ENGIN/STEP_A/cst[1] ), 
        .D(\MAIN/ENGIN/STEP_A/cst[3] ) );
    snl_invx05 \MAIN/ENGIN/STEP_A/deocgen_1/U13  ( .ZN(
        \MAIN/ENGIN/STEP_A/deocgen_1/n3543 ), .A(\MAIN/ENGIN/STEP_A/cst[2] )
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_B/deocgen_1/U12  ( .ZN(
        \MAIN/ENGIN/b_deocenh ), .A(\MAIN/ENGIN/STEP_B/cst[0] ), .B(
        \MAIN/ENGIN/STEP_B/deocgen_1/n3495 ), .C(\MAIN/ENGIN/STEP_B/cst[1] ), 
        .D(\MAIN/ENGIN/STEP_B/cst[3] ) );
    snl_invx05 \MAIN/ENGIN/STEP_B/deocgen_1/U13  ( .ZN(
        \MAIN/ENGIN/STEP_B/deocgen_1/n3495 ), .A(\MAIN/ENGIN/STEP_B/cst[2] )
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_C/deocgen_1/U12  ( .ZN(
        \MAIN/ENGIN/c_deocenh ), .A(\MAIN/ENGIN/STEP_C/cst[0] ), .B(
        \MAIN/ENGIN/STEP_C/deocgen_1/n3447 ), .C(\MAIN/ENGIN/STEP_C/cst[1] ), 
        .D(\MAIN/ENGIN/STEP_C/cst[3] ) );
    snl_invx05 \MAIN/ENGIN/STEP_C/deocgen_1/U13  ( .ZN(
        \MAIN/ENGIN/STEP_C/deocgen_1/n3447 ), .A(\MAIN/ENGIN/STEP_C/cst[2] )
         );
    snl_aoi112x0 \MAIN/ENGIN/STEP_D/deocgen_1/U12  ( .ZN(
        \MAIN/ENGIN/d_deocenh ), .A(\MAIN/ENGIN/STEP_D/cst[0] ), .B(
        \MAIN/ENGIN/STEP_D/deocgen_1/n3399 ), .C(\MAIN/ENGIN/STEP_D/cst[1] ), 
        .D(\MAIN/ENGIN/STEP_D/cst[3] ) );
    snl_invx05 \MAIN/ENGIN/STEP_D/deocgen_1/U13  ( .ZN(
        \MAIN/ENGIN/STEP_D/deocgen_1/n3399 ), .A(\MAIN/ENGIN/STEP_D/cst[2] )
         );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_7/U7  ( .Z(\ALUSHT/ALU/pkdecout[28] ), 
        .A(\ALUSHT/ALU/pkdecin[28] ), .B(\ALUSHT/ALU/dec32/gcarry[6] ), .C(
        \ALUSHT/ALU/dec32/dec4_7/n1796 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_7/U8  ( .Z(
        \ALUSHT/ALU/dec32/dec4_7/gg_out ), .A(\ALUSHT/ALU/pkdecin[28] ), .B(
        \ALUSHT/ALU/pkdecin[31] ), .C(\ALUSHT/ALU/pkdecin[29] ), .D(
        \ALUSHT/ALU/pkdecin[30] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_7/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_7/n1800 ), .A(\ALUSHT/ALU/dec32/dec4_7/n1796 ), 
        .B(\ALUSHT/ALU/dec32/dec4_7/n1799 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_7/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_7/n1798 ), .A(\ALUSHT/ALU/pkdecin[31] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_7/U9  ( .ZN(\ALUSHT/ALU/pkdecout[31] ), 
        .A(\ALUSHT/ALU/dec32/gcarry[6] ), .B(\ALUSHT/ALU/dec32/dec4_7/gg_out ), 
        .C(\ALUSHT/ALU/dec32/dec4_7/n1797 ), .D(
        \ALUSHT/ALU/dec32/dec4_7/n1798 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_7/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_7/n1796 ), .A(\ALUSHT/ALU/dec32/gcarry[6] ), 
        .B(\ALUSHT/ALU/pkdecin[28] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_7/U10  ( .ZN(\ALUSHT/ALU/pkdecout[29] 
        ), .A(\ALUSHT/ALU/dec32/dec4_7/n1796 ), .B(
        \ALUSHT/ALU/dec32/dec4_7/n1799 ), .C(\ALUSHT/ALU/dec32/dec4_7/n1800 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_7/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_7/n1799 ), .A(\ALUSHT/ALU/pkdecin[29] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_7/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_7/n1797 ), .A(\ALUSHT/ALU/pkdecin[30] ), .B(
        \ALUSHT/ALU/dec32/dec4_7/n1800 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_7/U16  ( .ZN(\ALUSHT/ALU/pkdecout[30] ), 
        .A(\ALUSHT/ALU/pkdecin[30] ), .B(\ALUSHT/ALU/dec32/dec4_7/n1800 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_0/U7  ( .Z(\ALUSHT/ALU/pkdecout[0] ), 
        .A(\ALUSHT/ALU/pkdecin[0] ), .B(1'b0), .C(
        \ALUSHT/ALU/dec32/dec4_0/n1791 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_0/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[0] ), 
        .A(\ALUSHT/ALU/pkdecin[0] ), .B(\ALUSHT/ALU/pkdecin[3] ), .C(
        \ALUSHT/ALU/pkdecin[1] ), .D(\ALUSHT/ALU/pkdecin[2] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_0/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_0/n1795 ), .A(\ALUSHT/ALU/dec32/dec4_0/n1791 ), 
        .B(\ALUSHT/ALU/dec32/dec4_0/n1794 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_0/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_0/n1793 ), .A(\ALUSHT/ALU/pkdecin[3] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_0/U9  ( .ZN(\ALUSHT/ALU/pkdecout[3] ), 
        .A(1'b0), .B(\ALUSHT/ALU/dec32/gg_out[0] ), .C(
        \ALUSHT/ALU/dec32/dec4_0/n1792 ), .D(\ALUSHT/ALU/dec32/dec4_0/n1793 )
         );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_0/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_0/n1791 ), .A(1'b0), .B(\ALUSHT/ALU/pkdecin[0] 
        ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_0/U10  ( .ZN(\ALUSHT/ALU/pkdecout[1] ), 
        .A(\ALUSHT/ALU/dec32/dec4_0/n1791 ), .B(
        \ALUSHT/ALU/dec32/dec4_0/n1794 ), .C(\ALUSHT/ALU/dec32/dec4_0/n1795 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_0/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_0/n1794 ), .A(\ALUSHT/ALU/pkdecin[1] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_0/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_0/n1792 ), .A(\ALUSHT/ALU/pkdecin[2] ), .B(
        \ALUSHT/ALU/dec32/dec4_0/n1795 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_0/U16  ( .ZN(\ALUSHT/ALU/pkdecout[2] ), 
        .A(\ALUSHT/ALU/pkdecin[2] ), .B(\ALUSHT/ALU/dec32/dec4_0/n1795 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_1/U7  ( .Z(\ALUSHT/ALU/pkdecout[4] ), 
        .A(\ALUSHT/ALU/pkdecin[4] ), .B(\ALUSHT/ALU/dec32/gg_out[0] ), .C(
        \ALUSHT/ALU/dec32/dec4_1/n1786 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_1/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[1] ), 
        .A(\ALUSHT/ALU/pkdecin[4] ), .B(\ALUSHT/ALU/pkdecin[7] ), .C(
        \ALUSHT/ALU/pkdecin[5] ), .D(\ALUSHT/ALU/pkdecin[6] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_1/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_1/n1790 ), .A(\ALUSHT/ALU/dec32/dec4_1/n1786 ), 
        .B(\ALUSHT/ALU/dec32/dec4_1/n1789 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_1/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_1/n1788 ), .A(\ALUSHT/ALU/pkdecin[7] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_1/U9  ( .ZN(\ALUSHT/ALU/pkdecout[7] ), 
        .A(\ALUSHT/ALU/dec32/gg_out[0] ), .B(\ALUSHT/ALU/dec32/gg_out[1] ), 
        .C(\ALUSHT/ALU/dec32/dec4_1/n1787 ), .D(
        \ALUSHT/ALU/dec32/dec4_1/n1788 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_1/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_1/n1786 ), .A(\ALUSHT/ALU/dec32/gg_out[0] ), 
        .B(\ALUSHT/ALU/pkdecin[4] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_1/U10  ( .ZN(\ALUSHT/ALU/pkdecout[5] ), 
        .A(\ALUSHT/ALU/dec32/dec4_1/n1786 ), .B(
        \ALUSHT/ALU/dec32/dec4_1/n1789 ), .C(\ALUSHT/ALU/dec32/dec4_1/n1790 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_1/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_1/n1789 ), .A(\ALUSHT/ALU/pkdecin[5] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_1/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_1/n1787 ), .A(\ALUSHT/ALU/pkdecin[6] ), .B(
        \ALUSHT/ALU/dec32/dec4_1/n1790 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_1/U16  ( .ZN(\ALUSHT/ALU/pkdecout[6] ), 
        .A(\ALUSHT/ALU/pkdecin[6] ), .B(\ALUSHT/ALU/dec32/dec4_1/n1790 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_2/U7  ( .Z(\ALUSHT/ALU/pkdecout[8] ), 
        .A(\ALUSHT/ALU/pkdecin[8] ), .B(\ALUSHT/ALU/dec32/gcarry[1] ), .C(
        \ALUSHT/ALU/dec32/dec4_2/n1781 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_2/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[2] ), 
        .A(\ALUSHT/ALU/pkdecin[8] ), .B(\ALUSHT/ALU/pkdecin[11] ), .C(
        \ALUSHT/ALU/pkdecin[9] ), .D(\ALUSHT/ALU/pkdecin[10] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_2/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_2/n1785 ), .A(\ALUSHT/ALU/dec32/dec4_2/n1781 ), 
        .B(\ALUSHT/ALU/dec32/dec4_2/n1784 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_2/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_2/n1783 ), .A(\ALUSHT/ALU/pkdecin[11] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_2/U9  ( .ZN(\ALUSHT/ALU/pkdecout[11] ), 
        .A(\ALUSHT/ALU/dec32/gcarry[1] ), .B(\ALUSHT/ALU/dec32/gg_out[2] ), 
        .C(\ALUSHT/ALU/dec32/dec4_2/n1782 ), .D(
        \ALUSHT/ALU/dec32/dec4_2/n1783 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_2/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_2/n1781 ), .A(\ALUSHT/ALU/dec32/gcarry[1] ), 
        .B(\ALUSHT/ALU/pkdecin[8] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_2/U10  ( .ZN(\ALUSHT/ALU/pkdecout[9] ), 
        .A(\ALUSHT/ALU/dec32/dec4_2/n1781 ), .B(
        \ALUSHT/ALU/dec32/dec4_2/n1784 ), .C(\ALUSHT/ALU/dec32/dec4_2/n1785 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_2/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_2/n1784 ), .A(\ALUSHT/ALU/pkdecin[9] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_2/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_2/n1782 ), .A(\ALUSHT/ALU/pkdecin[10] ), .B(
        \ALUSHT/ALU/dec32/dec4_2/n1785 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_2/U16  ( .ZN(\ALUSHT/ALU/pkdecout[10] ), 
        .A(\ALUSHT/ALU/pkdecin[10] ), .B(\ALUSHT/ALU/dec32/dec4_2/n1785 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_3/U7  ( .Z(\ALUSHT/ALU/pkdecout[12] ), 
        .A(\ALUSHT/ALU/pkdecin[12] ), .B(\ALUSHT/ALU/dec32/gcarry[2] ), .C(
        \ALUSHT/ALU/dec32/dec4_3/n1776 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_3/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[3] ), 
        .A(\ALUSHT/ALU/pkdecin[12] ), .B(\ALUSHT/ALU/pkdecin[15] ), .C(
        \ALUSHT/ALU/pkdecin[13] ), .D(\ALUSHT/ALU/pkdecin[14] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_3/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_3/n1780 ), .A(\ALUSHT/ALU/dec32/dec4_3/n1776 ), 
        .B(\ALUSHT/ALU/dec32/dec4_3/n1779 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_3/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_3/n1778 ), .A(\ALUSHT/ALU/pkdecin[15] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_3/U9  ( .ZN(\ALUSHT/ALU/pkdecout[15] ), 
        .A(\ALUSHT/ALU/dec32/gcarry[2] ), .B(\ALUSHT/ALU/dec32/gg_out[3] ), 
        .C(\ALUSHT/ALU/dec32/dec4_3/n1777 ), .D(
        \ALUSHT/ALU/dec32/dec4_3/n1778 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_3/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_3/n1776 ), .A(\ALUSHT/ALU/dec32/gcarry[2] ), 
        .B(\ALUSHT/ALU/pkdecin[12] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_3/U10  ( .ZN(\ALUSHT/ALU/pkdecout[13] 
        ), .A(\ALUSHT/ALU/dec32/dec4_3/n1776 ), .B(
        \ALUSHT/ALU/dec32/dec4_3/n1779 ), .C(\ALUSHT/ALU/dec32/dec4_3/n1780 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_3/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_3/n1779 ), .A(\ALUSHT/ALU/pkdecin[13] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_3/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_3/n1777 ), .A(\ALUSHT/ALU/pkdecin[14] ), .B(
        \ALUSHT/ALU/dec32/dec4_3/n1780 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_3/U16  ( .ZN(\ALUSHT/ALU/pkdecout[14] ), 
        .A(\ALUSHT/ALU/pkdecin[14] ), .B(\ALUSHT/ALU/dec32/dec4_3/n1780 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_4/U7  ( .Z(\ALUSHT/ALU/pkdecout[16] ), 
        .A(\ALUSHT/ALU/pkdecin[16] ), .B(\ALUSHT/ALU/dec32/gcarry[3] ), .C(
        \ALUSHT/ALU/dec32/dec4_4/n1771 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_4/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[4] ), 
        .A(\ALUSHT/ALU/pkdecin[16] ), .B(\ALUSHT/ALU/pkdecin[19] ), .C(
        \ALUSHT/ALU/pkdecin[17] ), .D(\ALUSHT/ALU/pkdecin[18] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_4/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_4/n1775 ), .A(\ALUSHT/ALU/dec32/dec4_4/n1771 ), 
        .B(\ALUSHT/ALU/dec32/dec4_4/n1774 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_4/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_4/n1773 ), .A(\ALUSHT/ALU/pkdecin[19] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_4/U9  ( .ZN(\ALUSHT/ALU/pkdecout[19] ), 
        .A(\ALUSHT/ALU/dec32/gcarry[3] ), .B(\ALUSHT/ALU/dec32/gg_out[4] ), 
        .C(\ALUSHT/ALU/dec32/dec4_4/n1772 ), .D(
        \ALUSHT/ALU/dec32/dec4_4/n1773 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_4/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_4/n1771 ), .A(\ALUSHT/ALU/dec32/gcarry[3] ), 
        .B(\ALUSHT/ALU/pkdecin[16] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_4/U10  ( .ZN(\ALUSHT/ALU/pkdecout[17] 
        ), .A(\ALUSHT/ALU/dec32/dec4_4/n1771 ), .B(
        \ALUSHT/ALU/dec32/dec4_4/n1774 ), .C(\ALUSHT/ALU/dec32/dec4_4/n1775 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_4/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_4/n1774 ), .A(\ALUSHT/ALU/pkdecin[17] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_4/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_4/n1772 ), .A(\ALUSHT/ALU/pkdecin[18] ), .B(
        \ALUSHT/ALU/dec32/dec4_4/n1775 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_4/U16  ( .ZN(\ALUSHT/ALU/pkdecout[18] ), 
        .A(\ALUSHT/ALU/pkdecin[18] ), .B(\ALUSHT/ALU/dec32/dec4_4/n1775 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_6/U7  ( .Z(\ALUSHT/ALU/pkdecout[24] ), 
        .A(\ALUSHT/ALU/pkdecin[24] ), .B(\ALUSHT/ALU/dec32/gcarry[5] ), .C(
        \ALUSHT/ALU/dec32/dec4_6/n1766 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_6/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[6] ), 
        .A(\ALUSHT/ALU/pkdecin[24] ), .B(\ALUSHT/ALU/pkdecin[27] ), .C(
        \ALUSHT/ALU/pkdecin[25] ), .D(\ALUSHT/ALU/pkdecin[26] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_6/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_6/n1770 ), .A(\ALUSHT/ALU/dec32/dec4_6/n1766 ), 
        .B(\ALUSHT/ALU/dec32/dec4_6/n1769 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_6/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_6/n1768 ), .A(\ALUSHT/ALU/pkdecin[27] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_6/U9  ( .ZN(\ALUSHT/ALU/pkdecout[27] ), 
        .A(\ALUSHT/ALU/dec32/gcarry[5] ), .B(\ALUSHT/ALU/dec32/gg_out[6] ), 
        .C(\ALUSHT/ALU/dec32/dec4_6/n1767 ), .D(
        \ALUSHT/ALU/dec32/dec4_6/n1768 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_6/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_6/n1766 ), .A(\ALUSHT/ALU/dec32/gcarry[5] ), 
        .B(\ALUSHT/ALU/pkdecin[24] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_6/U10  ( .ZN(\ALUSHT/ALU/pkdecout[25] 
        ), .A(\ALUSHT/ALU/dec32/dec4_6/n1766 ), .B(
        \ALUSHT/ALU/dec32/dec4_6/n1769 ), .C(\ALUSHT/ALU/dec32/dec4_6/n1770 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_6/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_6/n1769 ), .A(\ALUSHT/ALU/pkdecin[25] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_6/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_6/n1767 ), .A(\ALUSHT/ALU/pkdecin[26] ), .B(
        \ALUSHT/ALU/dec32/dec4_6/n1770 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_6/U16  ( .ZN(\ALUSHT/ALU/pkdecout[26] ), 
        .A(\ALUSHT/ALU/pkdecin[26] ), .B(\ALUSHT/ALU/dec32/dec4_6/n1770 ) );
    snl_ao012x1 \ALUSHT/ALU/dec32/dec4_5/U7  ( .Z(\ALUSHT/ALU/pkdecout[20] ), 
        .A(\ALUSHT/ALU/pkdecin[20] ), .B(\ALUSHT/ALU/dec32/gcarry[4] ), .C(
        \ALUSHT/ALU/dec32/dec4_5/n1636 ) );
    snl_or04x1 \ALUSHT/ALU/dec32/dec4_5/U8  ( .Z(\ALUSHT/ALU/dec32/gg_out[5] ), 
        .A(\ALUSHT/ALU/pkdecin[20] ), .B(\ALUSHT/ALU/pkdecin[23] ), .C(
        \ALUSHT/ALU/pkdecin[21] ), .D(\ALUSHT/ALU/pkdecin[22] ) );
    snl_nand02x1 \ALUSHT/ALU/dec32/dec4_5/U13  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_5/n1765 ), .A(\ALUSHT/ALU/dec32/dec4_5/n1636 ), 
        .B(\ALUSHT/ALU/dec32/dec4_5/n1764 ) );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_5/U14  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_5/n1763 ), .A(\ALUSHT/ALU/pkdecin[23] ) );
    snl_oai022x1 \ALUSHT/ALU/dec32/dec4_5/U9  ( .ZN(\ALUSHT/ALU/pkdecout[23] ), 
        .A(\ALUSHT/ALU/dec32/gcarry[4] ), .B(\ALUSHT/ALU/dec32/gg_out[5] ), 
        .C(\ALUSHT/ALU/dec32/dec4_5/n1637 ), .D(
        \ALUSHT/ALU/dec32/dec4_5/n1763 ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_5/U12  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_5/n1636 ), .A(\ALUSHT/ALU/dec32/gcarry[4] ), 
        .B(\ALUSHT/ALU/pkdecin[20] ) );
    snl_oai012x1 \ALUSHT/ALU/dec32/dec4_5/U10  ( .ZN(\ALUSHT/ALU/pkdecout[21] 
        ), .A(\ALUSHT/ALU/dec32/dec4_5/n1636 ), .B(
        \ALUSHT/ALU/dec32/dec4_5/n1764 ), .C(\ALUSHT/ALU/dec32/dec4_5/n1765 )
         );
    snl_invx05 \ALUSHT/ALU/dec32/dec4_5/U15  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_5/n1764 ), .A(\ALUSHT/ALU/pkdecin[21] ) );
    snl_nor02x1 \ALUSHT/ALU/dec32/dec4_5/U11  ( .ZN(
        \ALUSHT/ALU/dec32/dec4_5/n1637 ), .A(\ALUSHT/ALU/pkdecin[22] ), .B(
        \ALUSHT/ALU/dec32/dec4_5/n1765 ) );
    snl_xnor2x0 \ALUSHT/ALU/dec32/dec4_5/U16  ( .ZN(\ALUSHT/ALU/pkdecout[22] ), 
        .A(\ALUSHT/ALU/pkdecin[22] ), .B(\ALUSHT/ALU/dec32/dec4_5/n1765 ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add0/U7  ( .ZN(
        \ALUSHT/ALU/add32/add0/c_last ), .A(\ALUSHT/ALU/add32/add0/n1357 ), 
        .B(\ALUSHT/ALU/add32/add0/n1358 ), .C(\ALUSHT/ALU/add32/add0/n1359 )
         );
    snl_nor05x1 \ALUSHT/ALU/add32/add0/U8  ( .ZN(\ALUSHT/ALU/add32/gp_out[0] ), 
        .A(\ALUSHT/ALU/add32/add0/n1360 ), .B(\ALUSHT/ALU/add32/add0/n1357 ), 
        .C(\ALUSHT/ALU/add32/add0/n1361 ), .D(\ALUSHT/ALU/add32/add0/n1362 ), 
        .E(\ALUSHT/ALU/add32/add0/n1363 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U13  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1373 ), .A(\ALUSHT/ALU/add32/add0/n1372 ), .B(
        \ALUSHT/ALU/add32/add0/n1374 ) );
    snl_and12x1 \ALUSHT/ALU/add32/add0/U14  ( .Z(\ALUSHT/ALU/add32/add0/n1375 
        ), .A(\ALUSHT/ALU/add32/add0/n1360 ), .B(\ALUSHT/ALU/add32/add0/n1376 
        ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add0/U21  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1376 ), .A(\ALUSHT/ALU/pkaddina[0] ), .B(
        \ALUSHT/ALU/pkaddinb[0] ) );
    snl_invx05 \ALUSHT/ALU/add32/add0/U28  ( .ZN(\ALUSHT/ALU/add32/add0/n1378 
        ), .A(\ALUSHT/ALU/add32/add0/n1357 ) );
    snl_invx05 \ALUSHT/ALU/add32/add0/U33  ( .ZN(\ALUSHT/ALU/add32/add0/n1371 
        ), .A(\ALUSHT/ALU/add32/add0/n1374 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U34  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1360 ), .A(\ALUSHT/ALU/pkaddina[0] ), .B(
        \ALUSHT/ALU/pkaddinb[0] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add0/U41  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1359 ), .A(\ALUSHT/ALU/pkaddina[4] ), .B(
        \ALUSHT/ALU/pkaddinb[4] ) );
    snl_nand12x1 \ALUSHT/ALU/add32/add0/U46  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1381 ), .A(\ALUSHT/ALU/add32/add0/n1382 ), .B(
        \ALUSHT/ALU/add32/add0/n1386 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add0/U26  ( .Z(\ALUSHT/ALU/pkaddsum[0] ), .A(
        \ALUSHT/ALU/pkaddcin ), .B(\ALUSHT/ALU/add32/add0/n1375 ) );
    snl_ao01b2x0 \ALUSHT/ALU/add32/add0/U9  ( .Z(\ALUSHT/ALU/add32/gg_out[0] ), 
        .A(\ALUSHT/ALU/add32/add0/n1363 ), .B(\ALUSHT/ALU/add32/add0/n1364 ), 
        .C(\ALUSHT/ALU/add32/add0/n1365 ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add0/U12  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1369 ), .A(\ALUSHT/ALU/add32/add0/n1370 ), .B(
        \ALUSHT/ALU/add32/add0/n1371 ), .C(\ALUSHT/ALU/add32/add0/n1372 ) );
    snl_oai013x0 \ALUSHT/ALU/add32/add0/U35  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1380 ), .A(\ALUSHT/ALU/add32/add0/n1384 ), .B(
        \ALUSHT/ALU/add32/add0/n1360 ), .C(\ALUSHT/ALU/add32/add0/n1362 ), .D(
        \ALUSHT/ALU/add32/add0/n1385 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U27  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1357 ), .A(\ALUSHT/ALU/pkaddina[4] ), .B(
        \ALUSHT/ALU/pkaddinb[4] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add0/U40  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1358 ), .A(\ALUSHT/ALU/add32/add0/n1380 ), .B(
        \ALUSHT/ALU/add32/add0/n1387 ), .C(\ALUSHT/ALU/add32/add0/n1368 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add0/U20  ( .Z(\ALUSHT/ALU/pkaddsum[1] ), .A(
        \ALUSHT/ALU/add32/add0/n1370 ), .B(\ALUSHT/ALU/add32/add0/n1373 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U29  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1382 ), .A(\ALUSHT/ALU/pkaddina[2] ), .B(
        \ALUSHT/ALU/pkaddinb[2] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add0/U47  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1377 ), .A(\ALUSHT/ALU/add32/add0/n1385 ), .B(
        \ALUSHT/ALU/add32/add0/n1361 ), .C(\ALUSHT/ALU/add32/add0/n1388 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U10  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1366 ), .A(\ALUSHT/ALU/add32/add0/n1365 ), .B(
        \ALUSHT/ALU/add32/add0/n1363 ) );
    snl_aoi0b12x0 \ALUSHT/ALU/add32/add0/U15  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1364 ), .A(\ALUSHT/ALU/add32/add0/n1377 ), .B(
        \ALUSHT/ALU/add32/add0/n1378 ), .C(\ALUSHT/ALU/add32/add0/n1359 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add0/U17  ( .Z(\ALUSHT/ALU/pkaddsum[4] ), .A(
        \ALUSHT/ALU/add32/add0/n1379 ), .B(\ALUSHT/ALU/add32/add0/n1358 ) );
    snl_nand12x1 \ALUSHT/ALU/add32/add0/U22  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1362 ), .A(\ALUSHT/ALU/add32/add0/n1382 ), .B(
        \ALUSHT/ALU/add32/add0/n1371 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U32  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1374 ), .A(\ALUSHT/ALU/pkaddina[1] ), .B(
        \ALUSHT/ALU/pkaddinb[1] ) );
    snl_invx05 \ALUSHT/ALU/add32/add0/U39  ( .ZN(\ALUSHT/ALU/add32/add0/n1368 
        ), .A(\ALUSHT/ALU/add32/add0/n1388 ) );
    snl_invx05 \ALUSHT/ALU/add32/add0/U30  ( .ZN(\ALUSHT/ALU/add32/add0/n1372 
        ), .A(\ALUSHT/ALU/add32/add0/n1383 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U42  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1363 ), .A(\ALUSHT/ALU/pkaddina[5] ), .B(
        \ALUSHT/ALU/pkaddinb[5] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add0/U45  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1370 ), .A(\ALUSHT/ALU/add32/add0/n1360 ), .B(
        \ALUSHT/ALU/add32/add0/n1384 ), .C(\ALUSHT/ALU/add32/add0/n1376 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U11  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1367 ), .A(\ALUSHT/ALU/add32/add0/n1368 ), .B(
        \ALUSHT/ALU/add32/add0/n1361 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add0/U19  ( .Z(\ALUSHT/ALU/pkaddsum[2] ), .A(
        \ALUSHT/ALU/add32/add0/n1381 ), .B(\ALUSHT/ALU/add32/add0/n1369 ) );
    snl_oa122x1 \ALUSHT/ALU/add32/add0/U25  ( .Z(\ALUSHT/ALU/add32/add0/n1385 
        ), .A(\ALUSHT/ALU/add32/add0/n1376 ), .B(\ALUSHT/ALU/add32/add0/n1362 
        ), .C(\ALUSHT/ALU/add32/add0/n1382 ), .D(\ALUSHT/ALU/add32/add0/n1383 
        ), .E(\ALUSHT/ALU/add32/add0/n1386 ) );
    snl_invx05 \ALUSHT/ALU/add32/add0/U37  ( .ZN(\ALUSHT/ALU/add32/add0/n1387 
        ), .A(\ALUSHT/ALU/add32/add0/n1361 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add0/U16  ( .Z(\ALUSHT/ALU/pkaddsum[5] ), .A(
        \ALUSHT/ALU/add32/add0/c_last ), .B(\ALUSHT/ALU/add32/add0/n1366 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add0/U18  ( .Z(\ALUSHT/ALU/pkaddsum[3] ), .A(
        \ALUSHT/ALU/add32/add0/n1380 ), .B(\ALUSHT/ALU/add32/add0/n1367 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add0/U36  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1361 ), .A(\ALUSHT/ALU/pkaddina[3] ), .B(
        \ALUSHT/ALU/pkaddinb[3] ) );
    snl_and02x1 \ALUSHT/ALU/add32/add0/U43  ( .Z(\ALUSHT/ALU/add32/add0/n1365 
        ), .A(\ALUSHT/ALU/pkaddina[5] ), .B(\ALUSHT/ALU/pkaddinb[5] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add0/U23  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1383 ), .A(\ALUSHT/ALU/pkaddina[1] ), .B(
        \ALUSHT/ALU/pkaddinb[1] ) );
    snl_invx05 \ALUSHT/ALU/add32/add0/U24  ( .ZN(\ALUSHT/ALU/add32/add0/n1384 
        ), .A(\ALUSHT/ALU/pkaddcin ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add0/U31  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1386 ), .A(\ALUSHT/ALU/pkaddina[2] ), .B(
        \ALUSHT/ALU/pkaddinb[2] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add0/U38  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1388 ), .A(\ALUSHT/ALU/pkaddina[3] ), .B(
        \ALUSHT/ALU/pkaddinb[3] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add0/U44  ( .ZN(
        \ALUSHT/ALU/add32/add0/n1379 ), .A(\ALUSHT/ALU/add32/add0/n1378 ), .B(
        \ALUSHT/ALU/add32/add0/n1359 ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add1/U7  ( .ZN(
        \ALUSHT/ALU/add32/add1/c_last ), .A(\ALUSHT/ALU/add32/add1/n1325 ), 
        .B(\ALUSHT/ALU/add32/add1/n1326 ), .C(\ALUSHT/ALU/add32/add1/n1327 )
         );
    snl_nor05x1 \ALUSHT/ALU/add32/add1/U8  ( .ZN(\ALUSHT/ALU/add32/gp_out[1] ), 
        .A(\ALUSHT/ALU/add32/add1/n1328 ), .B(\ALUSHT/ALU/add32/add1/n1325 ), 
        .C(\ALUSHT/ALU/add32/add1/n1329 ), .D(\ALUSHT/ALU/add32/add1/n1330 ), 
        .E(\ALUSHT/ALU/add32/add1/n1331 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U13  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1341 ), .A(\ALUSHT/ALU/add32/add1/n1340 ), .B(
        \ALUSHT/ALU/add32/add1/n1342 ) );
    snl_and12x1 \ALUSHT/ALU/add32/add1/U14  ( .Z(\ALUSHT/ALU/add32/add1/n1343 
        ), .A(\ALUSHT/ALU/add32/add1/n1328 ), .B(\ALUSHT/ALU/add32/add1/n1344 
        ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add1/U21  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1344 ), .A(\ALUSHT/ALU/pkaddina[6] ), .B(
        \ALUSHT/ALU/pkaddinb[6] ) );
    snl_invx05 \ALUSHT/ALU/add32/add1/U28  ( .ZN(\ALUSHT/ALU/add32/add1/n1346 
        ), .A(\ALUSHT/ALU/add32/add1/n1325 ) );
    snl_invx05 \ALUSHT/ALU/add32/add1/U33  ( .ZN(\ALUSHT/ALU/add32/add1/n1339 
        ), .A(\ALUSHT/ALU/add32/add1/n1342 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U34  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1328 ), .A(\ALUSHT/ALU/pkaddina[6] ), .B(
        \ALUSHT/ALU/pkaddinb[6] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add1/U41  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1327 ), .A(\ALUSHT/ALU/pkaddina[10] ), .B(
        \ALUSHT/ALU/pkaddinb[10] ) );
    snl_nand12x1 \ALUSHT/ALU/add32/add1/U46  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1349 ), .A(\ALUSHT/ALU/add32/add1/n1350 ), .B(
        \ALUSHT/ALU/add32/add1/n1354 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add1/U26  ( .Z(\ALUSHT/ALU/pkaddsum[6] ), .A(
        \ALUSHT/ALU/add32/cin_stg[0] ), .B(\ALUSHT/ALU/add32/add1/n1343 ) );
    snl_ao01b2x0 \ALUSHT/ALU/add32/add1/U9  ( .Z(\ALUSHT/ALU/add32/gg_out[1] ), 
        .A(\ALUSHT/ALU/add32/add1/n1331 ), .B(\ALUSHT/ALU/add32/add1/n1332 ), 
        .C(\ALUSHT/ALU/add32/add1/n1333 ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add1/U12  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1337 ), .A(\ALUSHT/ALU/add32/add1/n1338 ), .B(
        \ALUSHT/ALU/add32/add1/n1339 ), .C(\ALUSHT/ALU/add32/add1/n1340 ) );
    snl_oai013x0 \ALUSHT/ALU/add32/add1/U35  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1348 ), .A(\ALUSHT/ALU/add32/add1/n1352 ), .B(
        \ALUSHT/ALU/add32/add1/n1328 ), .C(\ALUSHT/ALU/add32/add1/n1330 ), .D(
        \ALUSHT/ALU/add32/add1/n1353 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U27  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1325 ), .A(\ALUSHT/ALU/pkaddina[10] ), .B(
        \ALUSHT/ALU/pkaddinb[10] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add1/U40  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1326 ), .A(\ALUSHT/ALU/add32/add1/n1348 ), .B(
        \ALUSHT/ALU/add32/add1/n1355 ), .C(\ALUSHT/ALU/add32/add1/n1336 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add1/U20  ( .Z(\ALUSHT/ALU/pkaddsum[7] ), .A(
        \ALUSHT/ALU/add32/add1/n1338 ), .B(\ALUSHT/ALU/add32/add1/n1341 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U29  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1350 ), .A(\ALUSHT/ALU/pkaddina[8] ), .B(
        \ALUSHT/ALU/pkaddinb[8] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add1/U47  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1345 ), .A(\ALUSHT/ALU/add32/add1/n1353 ), .B(
        \ALUSHT/ALU/add32/add1/n1329 ), .C(\ALUSHT/ALU/add32/add1/n1356 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U10  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1334 ), .A(\ALUSHT/ALU/add32/add1/n1333 ), .B(
        \ALUSHT/ALU/add32/add1/n1331 ) );
    snl_aoi0b12x0 \ALUSHT/ALU/add32/add1/U15  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1332 ), .A(\ALUSHT/ALU/add32/add1/n1345 ), .B(
        \ALUSHT/ALU/add32/add1/n1346 ), .C(\ALUSHT/ALU/add32/add1/n1327 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add1/U17  ( .Z(\ALUSHT/ALU/pkaddsum[10] ), 
        .A(\ALUSHT/ALU/add32/add1/n1347 ), .B(\ALUSHT/ALU/add32/add1/n1326 )
         );
    snl_nand12x1 \ALUSHT/ALU/add32/add1/U22  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1330 ), .A(\ALUSHT/ALU/add32/add1/n1350 ), .B(
        \ALUSHT/ALU/add32/add1/n1339 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U32  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1342 ), .A(\ALUSHT/ALU/pkaddina[7] ), .B(
        \ALUSHT/ALU/pkaddinb[7] ) );
    snl_invx05 \ALUSHT/ALU/add32/add1/U39  ( .ZN(\ALUSHT/ALU/add32/add1/n1336 
        ), .A(\ALUSHT/ALU/add32/add1/n1356 ) );
    snl_invx05 \ALUSHT/ALU/add32/add1/U30  ( .ZN(\ALUSHT/ALU/add32/add1/n1340 
        ), .A(\ALUSHT/ALU/add32/add1/n1351 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U42  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1331 ), .A(\ALUSHT/ALU/pkaddina[11] ), .B(
        \ALUSHT/ALU/pkaddinb[11] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add1/U45  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1338 ), .A(\ALUSHT/ALU/add32/add1/n1328 ), .B(
        \ALUSHT/ALU/add32/add1/n1352 ), .C(\ALUSHT/ALU/add32/add1/n1344 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U11  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1335 ), .A(\ALUSHT/ALU/add32/add1/n1336 ), .B(
        \ALUSHT/ALU/add32/add1/n1329 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add1/U19  ( .Z(\ALUSHT/ALU/pkaddsum[8] ), .A(
        \ALUSHT/ALU/add32/add1/n1349 ), .B(\ALUSHT/ALU/add32/add1/n1337 ) );
    snl_oa122x1 \ALUSHT/ALU/add32/add1/U25  ( .Z(\ALUSHT/ALU/add32/add1/n1353 
        ), .A(\ALUSHT/ALU/add32/add1/n1344 ), .B(\ALUSHT/ALU/add32/add1/n1330 
        ), .C(\ALUSHT/ALU/add32/add1/n1350 ), .D(\ALUSHT/ALU/add32/add1/n1351 
        ), .E(\ALUSHT/ALU/add32/add1/n1354 ) );
    snl_invx05 \ALUSHT/ALU/add32/add1/U37  ( .ZN(\ALUSHT/ALU/add32/add1/n1355 
        ), .A(\ALUSHT/ALU/add32/add1/n1329 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add1/U16  ( .Z(\ALUSHT/ALU/pkaddsum[11] ), 
        .A(\ALUSHT/ALU/add32/add1/c_last ), .B(\ALUSHT/ALU/add32/add1/n1334 )
         );
    snl_xor2x0 \ALUSHT/ALU/add32/add1/U18  ( .Z(\ALUSHT/ALU/pkaddsum[9] ), .A(
        \ALUSHT/ALU/add32/add1/n1348 ), .B(\ALUSHT/ALU/add32/add1/n1335 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add1/U36  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1329 ), .A(\ALUSHT/ALU/pkaddina[9] ), .B(
        \ALUSHT/ALU/pkaddinb[9] ) );
    snl_and02x1 \ALUSHT/ALU/add32/add1/U43  ( .Z(\ALUSHT/ALU/add32/add1/n1333 
        ), .A(\ALUSHT/ALU/pkaddina[11] ), .B(\ALUSHT/ALU/pkaddinb[11] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add1/U23  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1351 ), .A(\ALUSHT/ALU/pkaddina[7] ), .B(
        \ALUSHT/ALU/pkaddinb[7] ) );
    snl_invx05 \ALUSHT/ALU/add32/add1/U24  ( .ZN(\ALUSHT/ALU/add32/add1/n1352 
        ), .A(\ALUSHT/ALU/add32/cin_stg[0] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add1/U31  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1354 ), .A(\ALUSHT/ALU/pkaddina[8] ), .B(
        \ALUSHT/ALU/pkaddinb[8] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add1/U38  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1356 ), .A(\ALUSHT/ALU/pkaddina[9] ), .B(
        \ALUSHT/ALU/pkaddinb[9] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add1/U44  ( .ZN(
        \ALUSHT/ALU/add32/add1/n1347 ), .A(\ALUSHT/ALU/add32/add1/n1346 ), .B(
        \ALUSHT/ALU/add32/add1/n1327 ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add2/U7  ( .ZN(
        \ALUSHT/ALU/add32/add2/c_last ), .A(\ALUSHT/ALU/add32/add2/n1293 ), 
        .B(\ALUSHT/ALU/add32/add2/n1294 ), .C(\ALUSHT/ALU/add32/add2/n1295 )
         );
    snl_nor05x1 \ALUSHT/ALU/add32/add2/U8  ( .ZN(\ALUSHT/ALU/add32/gp_out[2] ), 
        .A(\ALUSHT/ALU/add32/add2/n1296 ), .B(\ALUSHT/ALU/add32/add2/n1293 ), 
        .C(\ALUSHT/ALU/add32/add2/n1297 ), .D(\ALUSHT/ALU/add32/add2/n1298 ), 
        .E(\ALUSHT/ALU/add32/add2/n1299 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U13  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1309 ), .A(\ALUSHT/ALU/add32/add2/n1308 ), .B(
        \ALUSHT/ALU/add32/add2/n1310 ) );
    snl_and12x1 \ALUSHT/ALU/add32/add2/U14  ( .Z(\ALUSHT/ALU/add32/add2/n1311 
        ), .A(\ALUSHT/ALU/add32/add2/n1296 ), .B(\ALUSHT/ALU/add32/add2/n1312 
        ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add2/U21  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1312 ), .A(\ALUSHT/ALU/pkaddina[12] ), .B(
        \ALUSHT/ALU/pkaddinb[12] ) );
    snl_invx05 \ALUSHT/ALU/add32/add2/U28  ( .ZN(\ALUSHT/ALU/add32/add2/n1314 
        ), .A(\ALUSHT/ALU/add32/add2/n1293 ) );
    snl_invx05 \ALUSHT/ALU/add32/add2/U33  ( .ZN(\ALUSHT/ALU/add32/add2/n1307 
        ), .A(\ALUSHT/ALU/add32/add2/n1310 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U34  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1296 ), .A(\ALUSHT/ALU/pkaddina[12] ), .B(
        \ALUSHT/ALU/pkaddinb[12] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add2/U41  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1295 ), .A(\ALUSHT/ALU/pkaddina[16] ), .B(
        \ALUSHT/ALU/pkaddinb[16] ) );
    snl_nand12x1 \ALUSHT/ALU/add32/add2/U46  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1317 ), .A(\ALUSHT/ALU/add32/add2/n1318 ), .B(
        \ALUSHT/ALU/add32/add2/n1322 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add2/U26  ( .Z(\ALUSHT/ALU/pkaddsum[12] ), 
        .A(\ALUSHT/ALU/add32/cin_stg[1] ), .B(\ALUSHT/ALU/add32/add2/n1311 )
         );
    snl_ao01b2x0 \ALUSHT/ALU/add32/add2/U9  ( .Z(\ALUSHT/ALU/add32/gg_out[2] ), 
        .A(\ALUSHT/ALU/add32/add2/n1299 ), .B(\ALUSHT/ALU/add32/add2/n1300 ), 
        .C(\ALUSHT/ALU/add32/add2/n1301 ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add2/U12  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1305 ), .A(\ALUSHT/ALU/add32/add2/n1306 ), .B(
        \ALUSHT/ALU/add32/add2/n1307 ), .C(\ALUSHT/ALU/add32/add2/n1308 ) );
    snl_oai013x0 \ALUSHT/ALU/add32/add2/U35  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1316 ), .A(\ALUSHT/ALU/add32/add2/n1320 ), .B(
        \ALUSHT/ALU/add32/add2/n1296 ), .C(\ALUSHT/ALU/add32/add2/n1298 ), .D(
        \ALUSHT/ALU/add32/add2/n1321 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U27  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1293 ), .A(\ALUSHT/ALU/pkaddina[16] ), .B(
        \ALUSHT/ALU/pkaddinb[16] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add2/U40  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1294 ), .A(\ALUSHT/ALU/add32/add2/n1316 ), .B(
        \ALUSHT/ALU/add32/add2/n1323 ), .C(\ALUSHT/ALU/add32/add2/n1304 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add2/U20  ( .Z(\ALUSHT/ALU/pkaddsum[13] ), 
        .A(\ALUSHT/ALU/add32/add2/n1306 ), .B(\ALUSHT/ALU/add32/add2/n1309 )
         );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U29  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1318 ), .A(\ALUSHT/ALU/pkaddina[14] ), .B(
        \ALUSHT/ALU/pkaddinb[14] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add2/U47  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1313 ), .A(\ALUSHT/ALU/add32/add2/n1321 ), .B(
        \ALUSHT/ALU/add32/add2/n1297 ), .C(\ALUSHT/ALU/add32/add2/n1324 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U10  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1302 ), .A(\ALUSHT/ALU/add32/add2/n1301 ), .B(
        \ALUSHT/ALU/add32/add2/n1299 ) );
    snl_aoi0b12x0 \ALUSHT/ALU/add32/add2/U15  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1300 ), .A(\ALUSHT/ALU/add32/add2/n1313 ), .B(
        \ALUSHT/ALU/add32/add2/n1314 ), .C(\ALUSHT/ALU/add32/add2/n1295 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add2/U17  ( .Z(\ALUSHT/ALU/pkaddsum[16] ), 
        .A(\ALUSHT/ALU/add32/add2/n1315 ), .B(\ALUSHT/ALU/add32/add2/n1294 )
         );
    snl_nand12x1 \ALUSHT/ALU/add32/add2/U22  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1298 ), .A(\ALUSHT/ALU/add32/add2/n1318 ), .B(
        \ALUSHT/ALU/add32/add2/n1307 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U32  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1310 ), .A(\ALUSHT/ALU/pkaddina[13] ), .B(
        \ALUSHT/ALU/pkaddinb[13] ) );
    snl_invx05 \ALUSHT/ALU/add32/add2/U39  ( .ZN(\ALUSHT/ALU/add32/add2/n1304 
        ), .A(\ALUSHT/ALU/add32/add2/n1324 ) );
    snl_invx05 \ALUSHT/ALU/add32/add2/U30  ( .ZN(\ALUSHT/ALU/add32/add2/n1308 
        ), .A(\ALUSHT/ALU/add32/add2/n1319 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U42  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1299 ), .A(\ALUSHT/ALU/pkaddina[17] ), .B(
        \ALUSHT/ALU/pkaddinb[17] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add2/U45  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1306 ), .A(\ALUSHT/ALU/add32/add2/n1296 ), .B(
        \ALUSHT/ALU/add32/add2/n1320 ), .C(\ALUSHT/ALU/add32/add2/n1312 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U11  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1303 ), .A(\ALUSHT/ALU/add32/add2/n1304 ), .B(
        \ALUSHT/ALU/add32/add2/n1297 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add2/U19  ( .Z(\ALUSHT/ALU/pkaddsum[14] ), 
        .A(\ALUSHT/ALU/add32/add2/n1317 ), .B(\ALUSHT/ALU/add32/add2/n1305 )
         );
    snl_oa122x1 \ALUSHT/ALU/add32/add2/U25  ( .Z(\ALUSHT/ALU/add32/add2/n1321 
        ), .A(\ALUSHT/ALU/add32/add2/n1312 ), .B(\ALUSHT/ALU/add32/add2/n1298 
        ), .C(\ALUSHT/ALU/add32/add2/n1318 ), .D(\ALUSHT/ALU/add32/add2/n1319 
        ), .E(\ALUSHT/ALU/add32/add2/n1322 ) );
    snl_invx05 \ALUSHT/ALU/add32/add2/U37  ( .ZN(\ALUSHT/ALU/add32/add2/n1323 
        ), .A(\ALUSHT/ALU/add32/add2/n1297 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add2/U16  ( .Z(\ALUSHT/ALU/pkaddsum[17] ), 
        .A(\ALUSHT/ALU/add32/add2/c_last ), .B(\ALUSHT/ALU/add32/add2/n1302 )
         );
    snl_xor2x0 \ALUSHT/ALU/add32/add2/U18  ( .Z(\ALUSHT/ALU/pkaddsum[15] ), 
        .A(\ALUSHT/ALU/add32/add2/n1316 ), .B(\ALUSHT/ALU/add32/add2/n1303 )
         );
    snl_nor02x1 \ALUSHT/ALU/add32/add2/U36  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1297 ), .A(\ALUSHT/ALU/pkaddina[15] ), .B(
        \ALUSHT/ALU/pkaddinb[15] ) );
    snl_and02x1 \ALUSHT/ALU/add32/add2/U43  ( .Z(\ALUSHT/ALU/add32/add2/n1301 
        ), .A(\ALUSHT/ALU/pkaddina[17] ), .B(\ALUSHT/ALU/pkaddinb[17] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add2/U23  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1319 ), .A(\ALUSHT/ALU/pkaddina[13] ), .B(
        \ALUSHT/ALU/pkaddinb[13] ) );
    snl_invx05 \ALUSHT/ALU/add32/add2/U24  ( .ZN(\ALUSHT/ALU/add32/add2/n1320 
        ), .A(\ALUSHT/ALU/add32/cin_stg[1] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add2/U31  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1322 ), .A(\ALUSHT/ALU/pkaddina[14] ), .B(
        \ALUSHT/ALU/pkaddinb[14] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add2/U38  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1324 ), .A(\ALUSHT/ALU/pkaddina[15] ), .B(
        \ALUSHT/ALU/pkaddinb[15] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add2/U44  ( .ZN(
        \ALUSHT/ALU/add32/add2/n1315 ), .A(\ALUSHT/ALU/add32/add2/n1314 ), .B(
        \ALUSHT/ALU/add32/add2/n1295 ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add5/U7  ( .ZN(\ALUSHT/ALU/add32/c_last ), 
        .A(\ALUSHT/ALU/add32/add5/n1273 ), .B(\ALUSHT/ALU/add32/add5/n1274 ), 
        .C(\ALUSHT/ALU/add32/add5/n1275 ) );
    snl_nor04x0 \ALUSHT/ALU/add32/add5/U8  ( .ZN(\ALUSHT/ALU/add32/gp_out[5] ), 
        .A(\ALUSHT/ALU/add32/add5/n1273 ), .B(\ALUSHT/ALU/add32/add5/n1276 ), 
        .C(\ALUSHT/ALU/add32/add5/n1277 ), .D(\ALUSHT/ALU/add32/add5/n1278 )
         );
    snl_aoi0b12x0 \ALUSHT/ALU/add32/add5/U13  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1279 ), .A(\ALUSHT/ALU/add32/add5/n1286 ), .B(
        \ALUSHT/ALU/add32/add5/n1287 ), .C(\ALUSHT/ALU/add32/add5/n1275 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add5/U14  ( .Z(\ALUSHT/ALU/pkaddsum[31] ), 
        .A(\ALUSHT/ALU/add32/c_last ), .B(\ALUSHT/ALU/add32/add5/n1281 ) );
    snl_invx05 \ALUSHT/ALU/add32/add5/U21  ( .ZN(\ALUSHT/ALU/add32/add5/n1287 
        ), .A(\ALUSHT/ALU/add32/add5/n1273 ) );
    snl_aoi013x0 \ALUSHT/ALU/add32/add5/U28  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1274 ), .A(\ALUSHT/ALU/add32/cin_stg[4] ), .B(
        \ALUSHT/ALU/add32/add5/n1292 ), .C(\ALUSHT/ALU/add32/add5/n1283 ), .D(
        \ALUSHT/ALU/add32/add5/n1286 ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add5/U33  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1289 ), .A(\ALUSHT/ALU/add32/add5/n1292 ), .B(
        \ALUSHT/ALU/add32/add5/n1291 ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add5/U26  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1291 ), .A(\ALUSHT/ALU/pkaddina[29] ), .B(
        \ALUSHT/ALU/pkaddinb[29] ) );
    snl_ao01b2x0 \ALUSHT/ALU/add32/add5/U9  ( .Z(\ALUSHT/ALU/add32/gg_out[5] ), 
        .A(\ALUSHT/ALU/add32/add5/n1278 ), .B(\ALUSHT/ALU/add32/add5/n1279 ), 
        .C(\ALUSHT/ALU/add32/add5/n1280 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add5/U12  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1285 ), .A(\ALUSHT/ALU/add32/add5/n1284 ), .B(
        \ALUSHT/ALU/add32/add5/n1277 ) );
    snl_invx05 \ALUSHT/ALU/add32/add5/U27  ( .ZN(\ALUSHT/ALU/add32/add5/n1284 
        ), .A(\ALUSHT/ALU/add32/add5/n1290 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add5/U20  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1273 ), .A(\ALUSHT/ALU/pkaddina[30] ), .B(
        \ALUSHT/ALU/pkaddinb[30] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add5/U29  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1275 ), .A(\ALUSHT/ALU/pkaddina[30] ), .B(
        \ALUSHT/ALU/pkaddinb[30] ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add5/U10  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1281 ), .A(\ALUSHT/ALU/add32/add5/n1280 ), .B(
        \ALUSHT/ALU/add32/add5/n1278 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add5/U15  ( .Z(\ALUSHT/ALU/pkaddsum[30] ), 
        .A(\ALUSHT/ALU/add32/add5/n1288 ), .B(\ALUSHT/ALU/add32/add5/n1274 )
         );
    snl_nand02x1 \ALUSHT/ALU/add32/add5/U17  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1290 ), .A(\ALUSHT/ALU/pkaddina[28] ), .B(
        \ALUSHT/ALU/pkaddinb[28] ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add5/U22  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1276 ), .A(\ALUSHT/ALU/pkaddina[29] ), .B(
        \ALUSHT/ALU/pkaddinb[29] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add5/U32  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1288 ), .A(\ALUSHT/ALU/add32/add5/n1287 ), .B(
        \ALUSHT/ALU/add32/add5/n1275 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add5/U30  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1278 ), .A(\ALUSHT/ALU/pkaddina[31] ), .B(
        \ALUSHT/ALU/pkaddinb[31] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add5/U11  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1282 ), .A(\ALUSHT/ALU/add32/cin_stg[4] ), .B(
        \ALUSHT/ALU/add32/add5/n1283 ), .C(\ALUSHT/ALU/add32/add5/n1284 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add5/U19  ( .Z(\ALUSHT/ALU/pkaddsum[28] ), 
        .A(\ALUSHT/ALU/add32/cin_stg[4] ), .B(\ALUSHT/ALU/add32/add5/n1285 )
         );
    snl_invx05 \ALUSHT/ALU/add32/add5/U25  ( .ZN(\ALUSHT/ALU/add32/add5/n1283 
        ), .A(\ALUSHT/ALU/add32/add5/n1277 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add5/U16  ( .Z(\ALUSHT/ALU/pkaddsum[29] ), 
        .A(\ALUSHT/ALU/add32/add5/n1289 ), .B(\ALUSHT/ALU/add32/add5/n1282 )
         );
    snl_oai012x1 \ALUSHT/ALU/add32/add5/U18  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1286 ), .A(\ALUSHT/ALU/add32/add5/n1276 ), .B(
        \ALUSHT/ALU/add32/add5/n1290 ), .C(\ALUSHT/ALU/add32/add5/n1291 ) );
    snl_invx05 \ALUSHT/ALU/add32/add5/U23  ( .ZN(\ALUSHT/ALU/add32/add5/n1292 
        ), .A(\ALUSHT/ALU/add32/add5/n1276 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add5/U24  ( .ZN(
        \ALUSHT/ALU/add32/add5/n1277 ), .A(\ALUSHT/ALU/pkaddina[28] ), .B(
        \ALUSHT/ALU/pkaddinb[28] ) );
    snl_and02x1 \ALUSHT/ALU/add32/add5/U31  ( .Z(\ALUSHT/ALU/add32/add5/n1280 
        ), .A(\ALUSHT/ALU/pkaddina[31] ), .B(\ALUSHT/ALU/pkaddinb[31] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add3/U7  ( .ZN(
        \ALUSHT/ALU/add32/add3/c_last ), .A(\ALUSHT/ALU/add32/add3/n1241 ), 
        .B(\ALUSHT/ALU/add32/add3/n1242 ), .C(\ALUSHT/ALU/add32/add3/n1243 )
         );
    snl_nor05x1 \ALUSHT/ALU/add32/add3/U8  ( .ZN(\ALUSHT/ALU/add32/gp_out[3] ), 
        .A(\ALUSHT/ALU/add32/add3/n1244 ), .B(\ALUSHT/ALU/add32/add3/n1241 ), 
        .C(\ALUSHT/ALU/add32/add3/n1245 ), .D(\ALUSHT/ALU/add32/add3/n1246 ), 
        .E(\ALUSHT/ALU/add32/add3/n1247 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U13  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1257 ), .A(\ALUSHT/ALU/add32/add3/n1256 ), .B(
        \ALUSHT/ALU/add32/add3/n1258 ) );
    snl_and12x1 \ALUSHT/ALU/add32/add3/U14  ( .Z(\ALUSHT/ALU/add32/add3/n1259 
        ), .A(\ALUSHT/ALU/add32/add3/n1244 ), .B(\ALUSHT/ALU/add32/add3/n1260 
        ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add3/U21  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1260 ), .A(\ALUSHT/ALU/pkaddina[18] ), .B(
        \ALUSHT/ALU/pkaddinb[18] ) );
    snl_invx05 \ALUSHT/ALU/add32/add3/U28  ( .ZN(\ALUSHT/ALU/add32/add3/n1262 
        ), .A(\ALUSHT/ALU/add32/add3/n1241 ) );
    snl_invx05 \ALUSHT/ALU/add32/add3/U33  ( .ZN(\ALUSHT/ALU/add32/add3/n1255 
        ), .A(\ALUSHT/ALU/add32/add3/n1258 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U34  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1244 ), .A(\ALUSHT/ALU/pkaddina[18] ), .B(
        \ALUSHT/ALU/pkaddinb[18] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add3/U41  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1243 ), .A(\ALUSHT/ALU/pkaddina[22] ), .B(
        \ALUSHT/ALU/pkaddinb[22] ) );
    snl_nand12x1 \ALUSHT/ALU/add32/add3/U46  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1265 ), .A(\ALUSHT/ALU/add32/add3/n1266 ), .B(
        \ALUSHT/ALU/add32/add3/n1270 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add3/U26  ( .Z(\ALUSHT/ALU/pkaddsum[18] ), 
        .A(\ALUSHT/ALU/add32/cin_stg[2] ), .B(\ALUSHT/ALU/add32/add3/n1259 )
         );
    snl_ao01b2x0 \ALUSHT/ALU/add32/add3/U9  ( .Z(\ALUSHT/ALU/add32/gg_out[3] ), 
        .A(\ALUSHT/ALU/add32/add3/n1247 ), .B(\ALUSHT/ALU/add32/add3/n1248 ), 
        .C(\ALUSHT/ALU/add32/add3/n1249 ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add3/U12  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1253 ), .A(\ALUSHT/ALU/add32/add3/n1254 ), .B(
        \ALUSHT/ALU/add32/add3/n1255 ), .C(\ALUSHT/ALU/add32/add3/n1256 ) );
    snl_oai013x0 \ALUSHT/ALU/add32/add3/U35  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1264 ), .A(\ALUSHT/ALU/add32/add3/n1268 ), .B(
        \ALUSHT/ALU/add32/add3/n1244 ), .C(\ALUSHT/ALU/add32/add3/n1246 ), .D(
        \ALUSHT/ALU/add32/add3/n1269 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U27  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1241 ), .A(\ALUSHT/ALU/pkaddina[22] ), .B(
        \ALUSHT/ALU/pkaddinb[22] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add3/U40  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1242 ), .A(\ALUSHT/ALU/add32/add3/n1264 ), .B(
        \ALUSHT/ALU/add32/add3/n1271 ), .C(\ALUSHT/ALU/add32/add3/n1252 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add3/U20  ( .Z(\ALUSHT/ALU/pkaddsum[19] ), 
        .A(\ALUSHT/ALU/add32/add3/n1254 ), .B(\ALUSHT/ALU/add32/add3/n1257 )
         );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U29  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1266 ), .A(\ALUSHT/ALU/pkaddina[20] ), .B(
        \ALUSHT/ALU/pkaddinb[20] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add3/U47  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1261 ), .A(\ALUSHT/ALU/add32/add3/n1269 ), .B(
        \ALUSHT/ALU/add32/add3/n1245 ), .C(\ALUSHT/ALU/add32/add3/n1272 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U10  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1250 ), .A(\ALUSHT/ALU/add32/add3/n1249 ), .B(
        \ALUSHT/ALU/add32/add3/n1247 ) );
    snl_aoi0b12x0 \ALUSHT/ALU/add32/add3/U15  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1248 ), .A(\ALUSHT/ALU/add32/add3/n1261 ), .B(
        \ALUSHT/ALU/add32/add3/n1262 ), .C(\ALUSHT/ALU/add32/add3/n1243 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add3/U17  ( .Z(\ALUSHT/ALU/pkaddsum[22] ), 
        .A(\ALUSHT/ALU/add32/add3/n1263 ), .B(\ALUSHT/ALU/add32/add3/n1242 )
         );
    snl_nand12x1 \ALUSHT/ALU/add32/add3/U22  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1246 ), .A(\ALUSHT/ALU/add32/add3/n1266 ), .B(
        \ALUSHT/ALU/add32/add3/n1255 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U32  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1258 ), .A(\ALUSHT/ALU/pkaddina[19] ), .B(
        \ALUSHT/ALU/pkaddinb[19] ) );
    snl_invx05 \ALUSHT/ALU/add32/add3/U39  ( .ZN(\ALUSHT/ALU/add32/add3/n1252 
        ), .A(\ALUSHT/ALU/add32/add3/n1272 ) );
    snl_invx05 \ALUSHT/ALU/add32/add3/U30  ( .ZN(\ALUSHT/ALU/add32/add3/n1256 
        ), .A(\ALUSHT/ALU/add32/add3/n1267 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U42  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1247 ), .A(\ALUSHT/ALU/pkaddina[23] ), .B(
        \ALUSHT/ALU/pkaddinb[23] ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add3/U45  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1254 ), .A(\ALUSHT/ALU/add32/add3/n1244 ), .B(
        \ALUSHT/ALU/add32/add3/n1268 ), .C(\ALUSHT/ALU/add32/add3/n1260 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U11  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1251 ), .A(\ALUSHT/ALU/add32/add3/n1252 ), .B(
        \ALUSHT/ALU/add32/add3/n1245 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add3/U19  ( .Z(\ALUSHT/ALU/pkaddsum[20] ), 
        .A(\ALUSHT/ALU/add32/add3/n1265 ), .B(\ALUSHT/ALU/add32/add3/n1253 )
         );
    snl_oa122x1 \ALUSHT/ALU/add32/add3/U25  ( .Z(\ALUSHT/ALU/add32/add3/n1269 
        ), .A(\ALUSHT/ALU/add32/add3/n1260 ), .B(\ALUSHT/ALU/add32/add3/n1246 
        ), .C(\ALUSHT/ALU/add32/add3/n1266 ), .D(\ALUSHT/ALU/add32/add3/n1267 
        ), .E(\ALUSHT/ALU/add32/add3/n1270 ) );
    snl_invx05 \ALUSHT/ALU/add32/add3/U37  ( .ZN(\ALUSHT/ALU/add32/add3/n1271 
        ), .A(\ALUSHT/ALU/add32/add3/n1245 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add3/U16  ( .Z(\ALUSHT/ALU/pkaddsum[23] ), 
        .A(\ALUSHT/ALU/add32/add3/c_last ), .B(\ALUSHT/ALU/add32/add3/n1250 )
         );
    snl_xor2x0 \ALUSHT/ALU/add32/add3/U18  ( .Z(\ALUSHT/ALU/pkaddsum[21] ), 
        .A(\ALUSHT/ALU/add32/add3/n1264 ), .B(\ALUSHT/ALU/add32/add3/n1251 )
         );
    snl_nor02x1 \ALUSHT/ALU/add32/add3/U36  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1245 ), .A(\ALUSHT/ALU/pkaddina[21] ), .B(
        \ALUSHT/ALU/pkaddinb[21] ) );
    snl_and02x1 \ALUSHT/ALU/add32/add3/U43  ( .Z(\ALUSHT/ALU/add32/add3/n1249 
        ), .A(\ALUSHT/ALU/pkaddina[23] ), .B(\ALUSHT/ALU/pkaddinb[23] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add3/U23  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1267 ), .A(\ALUSHT/ALU/pkaddina[19] ), .B(
        \ALUSHT/ALU/pkaddinb[19] ) );
    snl_invx05 \ALUSHT/ALU/add32/add3/U24  ( .ZN(\ALUSHT/ALU/add32/add3/n1268 
        ), .A(\ALUSHT/ALU/add32/cin_stg[2] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add3/U31  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1270 ), .A(\ALUSHT/ALU/pkaddina[20] ), .B(
        \ALUSHT/ALU/pkaddinb[20] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add3/U38  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1272 ), .A(\ALUSHT/ALU/pkaddina[21] ), .B(
        \ALUSHT/ALU/pkaddinb[21] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add3/U44  ( .ZN(
        \ALUSHT/ALU/add32/add3/n1263 ), .A(\ALUSHT/ALU/add32/add3/n1262 ), .B(
        \ALUSHT/ALU/add32/add3/n1243 ) );
    snl_oai012x1 \ALUSHT/ALU/add32/add4/U7  ( .ZN(
        \ALUSHT/ALU/add32/add4/c_last ), .A(\ALUSHT/ALU/add32/add4/n1221 ), 
        .B(\ALUSHT/ALU/add32/add4/n1222 ), .C(\ALUSHT/ALU/add32/add4/n1223 )
         );
    snl_nor04x0 \ALUSHT/ALU/add32/add4/U8  ( .ZN(\ALUSHT/ALU/add32/gp_out[4] ), 
        .A(\ALUSHT/ALU/add32/add4/n1221 ), .B(\ALUSHT/ALU/add32/add4/n1224 ), 
        .C(\ALUSHT/ALU/add32/add4/n1225 ), .D(\ALUSHT/ALU/add32/add4/n1226 )
         );
    snl_aoi0b12x0 \ALUSHT/ALU/add32/add4/U13  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1227 ), .A(\ALUSHT/ALU/add32/add4/n1234 ), .B(
        \ALUSHT/ALU/add32/add4/n1235 ), .C(\ALUSHT/ALU/add32/add4/n1223 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add4/U14  ( .Z(\ALUSHT/ALU/pkaddsum[27] ), 
        .A(\ALUSHT/ALU/add32/add4/c_last ), .B(\ALUSHT/ALU/add32/add4/n1229 )
         );
    snl_invx05 \ALUSHT/ALU/add32/add4/U21  ( .ZN(\ALUSHT/ALU/add32/add4/n1235 
        ), .A(\ALUSHT/ALU/add32/add4/n1221 ) );
    snl_aoi013x0 \ALUSHT/ALU/add32/add4/U28  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1222 ), .A(\ALUSHT/ALU/add32/cin_stg[3] ), .B(
        \ALUSHT/ALU/add32/add4/n1240 ), .C(\ALUSHT/ALU/add32/add4/n1231 ), .D(
        \ALUSHT/ALU/add32/add4/n1234 ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add4/U33  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1237 ), .A(\ALUSHT/ALU/add32/add4/n1240 ), .B(
        \ALUSHT/ALU/add32/add4/n1239 ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add4/U26  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1239 ), .A(\ALUSHT/ALU/pkaddina[25] ), .B(
        \ALUSHT/ALU/pkaddinb[25] ) );
    snl_ao01b2x0 \ALUSHT/ALU/add32/add4/U9  ( .Z(\ALUSHT/ALU/add32/gg_out[4] ), 
        .A(\ALUSHT/ALU/add32/add4/n1226 ), .B(\ALUSHT/ALU/add32/add4/n1227 ), 
        .C(\ALUSHT/ALU/add32/add4/n1228 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add4/U12  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1233 ), .A(\ALUSHT/ALU/add32/add4/n1232 ), .B(
        \ALUSHT/ALU/add32/add4/n1225 ) );
    snl_invx05 \ALUSHT/ALU/add32/add4/U27  ( .ZN(\ALUSHT/ALU/add32/add4/n1232 
        ), .A(\ALUSHT/ALU/add32/add4/n1238 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add4/U20  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1221 ), .A(\ALUSHT/ALU/pkaddina[26] ), .B(
        \ALUSHT/ALU/pkaddinb[26] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add4/U29  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1223 ), .A(\ALUSHT/ALU/pkaddina[26] ), .B(
        \ALUSHT/ALU/pkaddinb[26] ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add4/U10  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1229 ), .A(\ALUSHT/ALU/add32/add4/n1228 ), .B(
        \ALUSHT/ALU/add32/add4/n1226 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add4/U15  ( .Z(\ALUSHT/ALU/pkaddsum[26] ), 
        .A(\ALUSHT/ALU/add32/add4/n1236 ), .B(\ALUSHT/ALU/add32/add4/n1222 )
         );
    snl_nand02x1 \ALUSHT/ALU/add32/add4/U17  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1238 ), .A(\ALUSHT/ALU/pkaddina[24] ), .B(
        \ALUSHT/ALU/pkaddinb[24] ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add4/U22  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1224 ), .A(\ALUSHT/ALU/pkaddina[25] ), .B(
        \ALUSHT/ALU/pkaddinb[25] ) );
    snl_nand02x1 \ALUSHT/ALU/add32/add4/U32  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1236 ), .A(\ALUSHT/ALU/add32/add4/n1235 ), .B(
        \ALUSHT/ALU/add32/add4/n1223 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add4/U30  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1226 ), .A(\ALUSHT/ALU/pkaddina[27] ), .B(
        \ALUSHT/ALU/pkaddinb[27] ) );
    snl_aoi012x1 \ALUSHT/ALU/add32/add4/U11  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1230 ), .A(\ALUSHT/ALU/add32/cin_stg[3] ), .B(
        \ALUSHT/ALU/add32/add4/n1231 ), .C(\ALUSHT/ALU/add32/add4/n1232 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add4/U19  ( .Z(\ALUSHT/ALU/pkaddsum[24] ), 
        .A(\ALUSHT/ALU/add32/cin_stg[3] ), .B(\ALUSHT/ALU/add32/add4/n1233 )
         );
    snl_invx05 \ALUSHT/ALU/add32/add4/U25  ( .ZN(\ALUSHT/ALU/add32/add4/n1231 
        ), .A(\ALUSHT/ALU/add32/add4/n1225 ) );
    snl_xor2x0 \ALUSHT/ALU/add32/add4/U16  ( .Z(\ALUSHT/ALU/pkaddsum[25] ), 
        .A(\ALUSHT/ALU/add32/add4/n1237 ), .B(\ALUSHT/ALU/add32/add4/n1230 )
         );
    snl_oai012x1 \ALUSHT/ALU/add32/add4/U18  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1234 ), .A(\ALUSHT/ALU/add32/add4/n1224 ), .B(
        \ALUSHT/ALU/add32/add4/n1238 ), .C(\ALUSHT/ALU/add32/add4/n1239 ) );
    snl_invx05 \ALUSHT/ALU/add32/add4/U23  ( .ZN(\ALUSHT/ALU/add32/add4/n1240 
        ), .A(\ALUSHT/ALU/add32/add4/n1224 ) );
    snl_nor02x1 \ALUSHT/ALU/add32/add4/U24  ( .ZN(
        \ALUSHT/ALU/add32/add4/n1225 ), .A(\ALUSHT/ALU/pkaddina[24] ), .B(
        \ALUSHT/ALU/pkaddinb[24] ) );
    snl_and02x1 \ALUSHT/ALU/add32/add4/U31  ( .Z(\ALUSHT/ALU/add32/add4/n1228 
        ), .A(\ALUSHT/ALU/pkaddina[27] ), .B(\ALUSHT/ALU/pkaddinb[27] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_7/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[7] ), .A(\ALUSHT/ALU/pkcmpinb[31] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_7/n1194 ), .C(\ALUSHT/ALU/cmp32/cmp4_7/n1195 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_7/n1196 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_7/U12  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_7/n1199 ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1200 ), 
        .B(\ALUSHT/ALU/intb[30] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_7/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_7/n1195 ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1194 ), 
        .B(\ALUSHT/ALU/pkcmpinb[31] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_7/U14  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[7] ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1201 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_7/n1202 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_7/n1203 ), .D(\ALUSHT/ALU/cmp32/cmp4_7/n1204 )
         );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1206 ), .A(\ALUSHT/ALU/intb[28] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1210 ), .A(\ALUSHT/ALU/pkcmpinb[31] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1208 ), .A(\ALUSHT/ALU/intb[30] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U15  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1205 ), .A(\ALUSHT/ALU/inta[29] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U20  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1196 ), .A(\ALUSHT/ALU/pkcmpina[31] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1209 ), .A(\ALUSHT/ALU/intb[29] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_7/U17  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_7/n1200 ), .A(\ALUSHT/ALU/intb[29] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_7/n1198 ), .C(\ALUSHT/ALU/cmp32/cmp4_7/n1197 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_7/n1205 ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_7/U22  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1201 ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1207 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_7/n1208 ), .C(\ALUSHT/ALU/inta[30] ), .D(
        \ALUSHT/ALU/intb[30] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_7/U11  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_7/n1197 ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1198 ), 
        .B(\ALUSHT/ALU/intb[29] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_7/U19  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_7/n1194 ), .A(\ALUSHT/ALU/intb[30] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_7/n1200 ), .C(\ALUSHT/ALU/cmp32/cmp4_7/n1199 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_7/n1207 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_7/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1202 ), .A(\ALUSHT/ALU/inta[28] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_7/n1206 ), .C(\ALUSHT/ALU/cmp32/cmp4_7/n1198 )
         );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_7/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1198 ), .A(\ALUSHT/ALU/inta[28] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_7/n1206 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_7/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1207 ), .A(\ALUSHT/ALU/inta[30] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_7/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1203 ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1205 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_7/n1209 ), .C(\ALUSHT/ALU/inta[29] ), .D(
        \ALUSHT/ALU/intb[29] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_7/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_7/n1204 ), .A(\ALUSHT/ALU/cmp32/cmp4_7/n1196 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_7/n1210 ), .C(\ALUSHT/ALU/pkcmpina[31] ), 
        .D(\ALUSHT/ALU/pkcmpinb[31] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_6/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[6] ), .A(\ALUSHT/ALU/intb[27] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_6/n1177 ), .C(\ALUSHT/ALU/cmp32/cmp4_6/n1178 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_6/n1179 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_6/U12  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_6/n1182 ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1183 ), 
        .B(\ALUSHT/ALU/intb[26] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_6/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_6/n1178 ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1177 ), 
        .B(\ALUSHT/ALU/intb[27] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_6/U14  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[6] ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1184 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_6/n1185 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_6/n1186 ), .D(\ALUSHT/ALU/cmp32/cmp4_6/n1187 )
         );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1189 ), .A(\ALUSHT/ALU/intb[24] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1193 ), .A(\ALUSHT/ALU/intb[27] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1191 ), .A(\ALUSHT/ALU/intb[26] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U15  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1188 ), .A(\ALUSHT/ALU/inta[25] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U20  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1179 ), .A(\ALUSHT/ALU/inta[27] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1192 ), .A(\ALUSHT/ALU/intb[25] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_6/U17  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_6/n1183 ), .A(\ALUSHT/ALU/intb[25] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_6/n1181 ), .C(\ALUSHT/ALU/cmp32/cmp4_6/n1180 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_6/n1188 ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_6/U22  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1184 ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1190 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_6/n1191 ), .C(\ALUSHT/ALU/inta[26] ), .D(
        \ALUSHT/ALU/intb[26] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_6/U11  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_6/n1180 ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1181 ), 
        .B(\ALUSHT/ALU/intb[25] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_6/U19  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_6/n1177 ), .A(\ALUSHT/ALU/intb[26] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_6/n1183 ), .C(\ALUSHT/ALU/cmp32/cmp4_6/n1182 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_6/n1190 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_6/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1185 ), .A(\ALUSHT/ALU/inta[24] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_6/n1189 ), .C(\ALUSHT/ALU/cmp32/cmp4_6/n1181 )
         );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_6/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1181 ), .A(\ALUSHT/ALU/inta[24] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_6/n1189 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_6/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1190 ), .A(\ALUSHT/ALU/inta[26] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_6/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1186 ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1188 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_6/n1192 ), .C(\ALUSHT/ALU/inta[25] ), .D(
        \ALUSHT/ALU/intb[25] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_6/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_6/n1187 ), .A(\ALUSHT/ALU/cmp32/cmp4_6/n1179 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_6/n1193 ), .C(\ALUSHT/ALU/inta[27] ), .D(
        \ALUSHT/ALU/intb[27] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_1/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1169 ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1171 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_1/n1175 ), .C(\pgaluina[5] ), .D(
        \pgaluinb[5] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_1/U12  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[1] ), .A(\pgaluinb[7] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_1/n1160 ), .C(\ALUSHT/ALU/cmp32/cmp4_1/n1161 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_1/n1162 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_1/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_1/n1163 ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1164 ), 
        .B(\pgaluinb[5] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_1/U14  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_1/n1165 ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1166 ), 
        .B(\pgaluinb[6] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_1/U21  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_1/n1160 ), .A(\pgaluinb[6] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_1/n1166 ), .C(\ALUSHT/ALU/cmp32/cmp4_1/n1165 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_1/n1173 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1176 ), .A(\pgaluinb[7] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1174 ), .A(\pgaluinb[6] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_1/U15  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_1/n1161 ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1160 ), 
        .B(\pgaluinb[7] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U20  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1173 ), .A(\pgaluina[6] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1175 ), .A(\pgaluinb[5] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U17  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1171 ), .A(\pgaluina[5] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U22  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1162 ), .A(\pgaluina[7] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_1/U11  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1170 ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1162 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_1/n1176 ), .C(\pgaluina[7] ), .D(
        \pgaluinb[7] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_1/U19  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_1/n1166 ), .A(\pgaluinb[5] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_1/n1164 ), .C(\ALUSHT/ALU/cmp32/cmp4_1/n1163 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_1/n1171 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_1/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1168 ), .A(\pgaluina[4] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_1/n1172 ), .C(\ALUSHT/ALU/cmp32/cmp4_1/n1164 )
         );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_1/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[1] ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1167 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_1/n1168 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_1/n1169 ), .D(\ALUSHT/ALU/cmp32/cmp4_1/n1170 )
         );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_1/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1164 ), .A(\pgaluina[4] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_1/n1172 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_1/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1172 ), .A(\pgaluinb[4] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_1/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_1/n1167 ), .A(\ALUSHT/ALU/cmp32/cmp4_1/n1173 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_1/n1174 ), .C(\pgaluina[6] ), .D(
        \pgaluinb[6] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_0/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1150 ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1156 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_0/n1157 ), .C(\pgaluina[2] ), .D(
        \pgaluinb[2] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_0/U12  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1153 ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1145 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_0/n1159 ), .C(\pgaluina[3] ), .D(
        \pgaluinb[3] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_0/U13  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[0] ), .A(\pgaluinb[3] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_0/n1143 ), .C(\ALUSHT/ALU/cmp32/cmp4_0/n1144 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_0/n1145 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_0/U14  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_0/n1146 ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1147 ), 
        .B(\pgaluinb[1] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1156 ), .A(\pgaluina[2] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1159 ), .A(\pgaluinb[3] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1157 ), .A(\pgaluinb[2] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_0/U15  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_0/n1148 ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1149 ), 
        .B(\pgaluinb[2] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_0/U20  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_0/n1149 ), .A(\pgaluinb[1] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_0/n1147 ), .C(\ALUSHT/ALU/cmp32/cmp4_0/n1146 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_0/n1154 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1158 ), .A(\pgaluinb[1] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_0/U17  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[0] ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1150 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_0/n1151 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_0/n1152 ), .D(\ALUSHT/ALU/cmp32/cmp4_0/n1153 )
         );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_0/U22  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_0/n1143 ), .A(\pgaluinb[2] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_0/n1149 ), .C(\ALUSHT/ALU/cmp32/cmp4_0/n1148 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_0/n1156 ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_0/U11  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1152 ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1154 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_0/n1158 ), .C(\pgaluina[1] ), .D(
        \pgaluinb[1] ) );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_0/U19  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1147 ), .A(\pgaluina[0] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_0/n1155 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_0/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1151 ), .A(\pgaluina[0] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_0/n1155 ), .C(\ALUSHT/ALU/cmp32/cmp4_0/n1147 )
         );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_0/U16  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_0/n1144 ), .A(\ALUSHT/ALU/cmp32/cmp4_0/n1143 ), 
        .B(\pgaluinb[3] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1154 ), .A(\pgaluina[1] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1145 ), .A(\pgaluina[3] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_0/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_0/n1155 ), .A(\pgaluinb[0] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_5/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[5] ), .A(\ALUSHT/ALU/intb[23] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_5/n1126 ), .C(\ALUSHT/ALU/cmp32/cmp4_5/n1127 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_5/n1128 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_5/U12  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_5/n1131 ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1132 ), 
        .B(\ALUSHT/ALU/intb[22] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_5/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_5/n1127 ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1126 ), 
        .B(\ALUSHT/ALU/intb[23] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_5/U14  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[5] ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1133 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_5/n1134 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_5/n1135 ), .D(\ALUSHT/ALU/cmp32/cmp4_5/n1136 )
         );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1138 ), .A(\ALUSHT/ALU/intb[20] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1142 ), .A(\ALUSHT/ALU/intb[23] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1140 ), .A(\ALUSHT/ALU/intb[22] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U15  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1137 ), .A(\ALUSHT/ALU/inta[21] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U20  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1128 ), .A(\ALUSHT/ALU/inta[23] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1141 ), .A(\ALUSHT/ALU/intb[21] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_5/U17  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_5/n1132 ), .A(\ALUSHT/ALU/intb[21] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_5/n1130 ), .C(\ALUSHT/ALU/cmp32/cmp4_5/n1129 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_5/n1137 ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_5/U22  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1133 ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1139 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_5/n1140 ), .C(\ALUSHT/ALU/inta[22] ), .D(
        \ALUSHT/ALU/intb[22] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_5/U11  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_5/n1129 ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1130 ), 
        .B(\ALUSHT/ALU/intb[21] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_5/U19  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_5/n1126 ), .A(\ALUSHT/ALU/intb[22] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_5/n1132 ), .C(\ALUSHT/ALU/cmp32/cmp4_5/n1131 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_5/n1139 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_5/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1134 ), .A(\ALUSHT/ALU/inta[20] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_5/n1138 ), .C(\ALUSHT/ALU/cmp32/cmp4_5/n1130 )
         );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_5/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1130 ), .A(\ALUSHT/ALU/inta[20] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_5/n1138 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_5/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1139 ), .A(\ALUSHT/ALU/inta[22] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_5/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1135 ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1137 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_5/n1141 ), .C(\ALUSHT/ALU/inta[21] ), .D(
        \ALUSHT/ALU/intb[21] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_5/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_5/n1136 ), .A(\ALUSHT/ALU/cmp32/cmp4_5/n1128 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_5/n1142 ), .C(\ALUSHT/ALU/inta[23] ), .D(
        \ALUSHT/ALU/intb[23] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_4/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[4] ), .A(\ALUSHT/ALU/intb[19] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_4/n1109 ), .C(\ALUSHT/ALU/cmp32/cmp4_4/n1110 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_4/n1111 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_4/U12  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_4/n1114 ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1115 ), 
        .B(\ALUSHT/ALU/intb[18] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_4/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_4/n1110 ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1109 ), 
        .B(\ALUSHT/ALU/intb[19] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_4/U14  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[4] ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1116 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_4/n1117 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_4/n1118 ), .D(\ALUSHT/ALU/cmp32/cmp4_4/n1119 )
         );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1121 ), .A(\ALUSHT/ALU/intb[16] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1125 ), .A(\ALUSHT/ALU/intb[19] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1123 ), .A(\ALUSHT/ALU/intb[18] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U15  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1120 ), .A(\ALUSHT/ALU/inta[17] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U20  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1111 ), .A(\ALUSHT/ALU/inta[19] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1124 ), .A(\ALUSHT/ALU/intb[17] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_4/U17  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_4/n1115 ), .A(\ALUSHT/ALU/intb[17] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_4/n1113 ), .C(\ALUSHT/ALU/cmp32/cmp4_4/n1112 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_4/n1120 ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_4/U22  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1116 ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1122 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_4/n1123 ), .C(\ALUSHT/ALU/inta[18] ), .D(
        \ALUSHT/ALU/intb[18] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_4/U11  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_4/n1112 ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1113 ), 
        .B(\ALUSHT/ALU/intb[17] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_4/U19  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_4/n1109 ), .A(\ALUSHT/ALU/intb[18] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_4/n1115 ), .C(\ALUSHT/ALU/cmp32/cmp4_4/n1114 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_4/n1122 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_4/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1117 ), .A(\ALUSHT/ALU/inta[16] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_4/n1121 ), .C(\ALUSHT/ALU/cmp32/cmp4_4/n1113 )
         );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_4/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1113 ), .A(\ALUSHT/ALU/inta[16] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_4/n1121 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_4/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1122 ), .A(\ALUSHT/ALU/inta[18] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_4/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1118 ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1120 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_4/n1124 ), .C(\ALUSHT/ALU/inta[17] ), .D(
        \ALUSHT/ALU/intb[17] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_4/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_4/n1119 ), .A(\ALUSHT/ALU/cmp32/cmp4_4/n1111 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_4/n1125 ), .C(\ALUSHT/ALU/inta[19] ), .D(
        \ALUSHT/ALU/intb[19] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_3/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1099 ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1105 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_3/n1106 ), .C(\pgaluina[14] ), .D(
        \pgaluinb[14] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_3/U12  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_3/n1095 ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1096 ), 
        .B(\pgaluinb[13] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_3/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_3/n1097 ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1098 ), 
        .B(\pgaluinb[14] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_3/U14  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_3/n1093 ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1092 ), 
        .B(\pgaluinb[15] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1094 ), .A(\pgaluina[15] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U28  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1108 ), .A(\pgaluinb[15] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U26  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1106 ), .A(\pgaluinb[14] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_3/U15  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[3] ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1099 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_3/n1100 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_3/n1101 ), .D(\ALUSHT/ALU/cmp32/cmp4_3/n1102 )
         );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_3/U20  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_3/n1092 ), .A(\pgaluinb[14] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_3/n1098 ), .C(\ALUSHT/ALU/cmp32/cmp4_3/n1097 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_3/n1105 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U27  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1107 ), .A(\pgaluinb[13] ) );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_3/U17  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1096 ), .A(\pgaluina[12] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_3/n1104 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U22  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1104 ), .A(\pgaluinb[12] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_3/U11  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[3] ), .A(\pgaluinb[15] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_3/n1092 ), .C(\ALUSHT/ALU/cmp32/cmp4_3/n1093 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_3/n1094 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U19  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1105 ), .A(\pgaluina[14] ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_3/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1100 ), .A(\pgaluina[12] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_3/n1104 ), .C(\ALUSHT/ALU/cmp32/cmp4_3/n1096 )
         );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_3/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1103 ), .A(\pgaluina[13] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_3/U18  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_3/n1098 ), .A(\pgaluinb[13] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_3/n1096 ), .C(\ALUSHT/ALU/cmp32/cmp4_3/n1095 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_3/n1103 ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_3/U23  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1101 ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1103 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_3/n1107 ), .C(\pgaluina[13] ), .D(
        \pgaluinb[13] ) );
    snl_aoi022x1 \ALUSHT/ALU/cmp32/cmp4_3/U24  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_3/n1102 ), .A(\ALUSHT/ALU/cmp32/cmp4_3/n1094 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_3/n1108 ), .C(\pgaluina[15] ), .D(
        \pgaluinb[15] ) );
    snl_oai022x1 \ALUSHT/ALU/cmp32/cmp4_2/U10  ( .ZN(
        \ALUSHT/ALU/cmp32/ggflg[2] ), .A(\pgaluinb[11] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_2/n1078 ), .C(\ALUSHT/ALU/cmp32/cmp4_2/n1079 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_2/n1080 ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_2/U12  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1083 ), .A(\ALUSHT/ALU/cmp32/cmp4_2/n1084 ), 
        .B(\pgaluinb[10] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_2/U13  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1079 ), .A(\ALUSHT/ALU/cmp32/cmp4_2/n1078 ), 
        .B(\pgaluinb[11] ) );
    snl_nor04x0 \ALUSHT/ALU/cmp32/cmp4_2/U14  ( .ZN(
        \ALUSHT/ALU/cmp32/geqflg[2] ), .A(\ALUSHT/ALU/cmp32/cmp4_2/n1085 ), 
        .B(\ALUSHT/ALU/cmp32/cmp4_2/n1086 ), .C(
        \ALUSHT/ALU/cmp32/cmp4_2/n1087 ), .D(\ALUSHT/ALU/cmp32/cmp4_2/n1088 )
         );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_2/U21  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_2/n1090 ), .A(\pgaluinb[8] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_2/U15  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_2/n1089 ), .A(\pgaluina[9] ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_2/U20  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_2/n1080 ), .A(\pgaluina[11] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_2/U17  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1084 ), .A(\pgaluinb[9] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_2/n1082 ), .C(\ALUSHT/ALU/cmp32/cmp4_2/n1081 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_2/n1089 ) );
    snl_xor2x0 \ALUSHT/ALU/cmp32/cmp4_2/U22  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1085 ), .A(\pgaluina[10] ), .B(
        \pgaluinb[10] ) );
    snl_and02x1 \ALUSHT/ALU/cmp32/cmp4_2/U11  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1081 ), .A(\ALUSHT/ALU/cmp32/cmp4_2/n1082 ), 
        .B(\pgaluinb[9] ) );
    snl_oa022x1 \ALUSHT/ALU/cmp32/cmp4_2/U19  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1078 ), .A(\pgaluinb[10] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_2/n1084 ), .C(\ALUSHT/ALU/cmp32/cmp4_2/n1083 ), 
        .D(\ALUSHT/ALU/cmp32/cmp4_2/n1091 ) );
    snl_oai012x1 \ALUSHT/ALU/cmp32/cmp4_2/U25  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_2/n1086 ), .A(\pgaluina[8] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_2/n1090 ), .C(\ALUSHT/ALU/cmp32/cmp4_2/n1082 )
         );
    snl_nand02x1 \ALUSHT/ALU/cmp32/cmp4_2/U16  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_2/n1082 ), .A(\pgaluina[8] ), .B(
        \ALUSHT/ALU/cmp32/cmp4_2/n1090 ) );
    snl_invx05 \ALUSHT/ALU/cmp32/cmp4_2/U18  ( .ZN(
        \ALUSHT/ALU/cmp32/cmp4_2/n1091 ), .A(\pgaluina[10] ) );
    snl_xor2x0 \ALUSHT/ALU/cmp32/cmp4_2/U23  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1087 ), .A(\pgaluina[9] ), .B(\pgaluinb[9] )
         );
    snl_xor2x0 \ALUSHT/ALU/cmp32/cmp4_2/U24  ( .Z(
        \ALUSHT/ALU/cmp32/cmp4_2/n1088 ), .A(\pgaluina[11] ), .B(
        \pgaluinb[11] ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_0/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[0] 
        ), .A(\ALUSHT/ALU/pkincin[3] ), .B(\ALUSHT/ALU/pkincin[0] ), .C(
        \ALUSHT/ALU/pkincin[1] ), .D(\ALUSHT/ALU/pkincin[2] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_0/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_0/n1075 ), .A(\ALUSHT/ALU/pkincin[0] ), .B(1'b1
        ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_0/U13  ( .Z(\ALUSHT/ALU/pkincout[0] ), 
        .A(\ALUSHT/ALU/pkincin[0] ), .B(1'b1) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_0/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_0/n1077 ), .A(\ALUSHT/ALU/pkincin[2] ), .B(
        \ALUSHT/ALU/inc32/inc4_0/n1076 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_0/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_0/n1076 ), .A(\ALUSHT/ALU/inc32/inc4_0/n1075 ), 
        .B(\ALUSHT/ALU/pkincin[1] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_0/U12  ( .ZN(\ALUSHT/ALU/pkincout[1] ), 
        .A(\ALUSHT/ALU/pkincin[1] ), .B(\ALUSHT/ALU/inc32/inc4_0/n1075 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_0/U10  ( .ZN(\ALUSHT/ALU/pkincout[3] ), 
        .A(\ALUSHT/ALU/pkincin[3] ), .B(\ALUSHT/ALU/inc32/inc4_0/n1077 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_0/U11  ( .Z(\ALUSHT/ALU/pkincout[2] ), 
        .A(\ALUSHT/ALU/pkincin[2] ), .B(\ALUSHT/ALU/inc32/inc4_0/n1076 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_1/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[1] 
        ), .A(\ALUSHT/ALU/pkincin[7] ), .B(\ALUSHT/ALU/pkincin[4] ), .C(
        \ALUSHT/ALU/pkincin[5] ), .D(\ALUSHT/ALU/pkincin[6] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_1/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_1/n1072 ), .A(\ALUSHT/ALU/pkincin[4] ), .B(
        \ALUSHT/ALU/inc32/gp_out[0] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_1/U13  ( .Z(\ALUSHT/ALU/pkincout[4] ), 
        .A(\ALUSHT/ALU/pkincin[4] ), .B(\ALUSHT/ALU/inc32/gp_out[0] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_1/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_1/n1074 ), .A(\ALUSHT/ALU/pkincin[6] ), .B(
        \ALUSHT/ALU/inc32/inc4_1/n1073 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_1/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_1/n1073 ), .A(\ALUSHT/ALU/inc32/inc4_1/n1072 ), 
        .B(\ALUSHT/ALU/pkincin[5] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_1/U12  ( .ZN(\ALUSHT/ALU/pkincout[5] ), 
        .A(\ALUSHT/ALU/pkincin[5] ), .B(\ALUSHT/ALU/inc32/inc4_1/n1072 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_1/U10  ( .ZN(\ALUSHT/ALU/pkincout[7] ), 
        .A(\ALUSHT/ALU/pkincin[7] ), .B(\ALUSHT/ALU/inc32/inc4_1/n1074 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_1/U11  ( .Z(\ALUSHT/ALU/pkincout[6] ), 
        .A(\ALUSHT/ALU/pkincin[6] ), .B(\ALUSHT/ALU/inc32/inc4_1/n1073 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_6/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[6] 
        ), .A(\ALUSHT/ALU/pkincin[27] ), .B(\ALUSHT/ALU/pkincin[24] ), .C(
        \ALUSHT/ALU/pkincin[25] ), .D(\ALUSHT/ALU/pkincin[26] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_6/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_6/n1069 ), .A(\ALUSHT/ALU/pkincin[24] ), .B(
        \ALUSHT/ALU/inc32/gg_out[5] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_6/U13  ( .Z(\ALUSHT/ALU/pkincout[24] ), 
        .A(\ALUSHT/ALU/pkincin[24] ), .B(\ALUSHT/ALU/inc32/gg_out[5] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_6/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_6/n1071 ), .A(\ALUSHT/ALU/pkincin[26] ), .B(
        \ALUSHT/ALU/inc32/inc4_6/n1070 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_6/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_6/n1070 ), .A(\ALUSHT/ALU/inc32/inc4_6/n1069 ), 
        .B(\ALUSHT/ALU/pkincin[25] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_6/U12  ( .ZN(\ALUSHT/ALU/pkincout[25] ), 
        .A(\ALUSHT/ALU/pkincin[25] ), .B(\ALUSHT/ALU/inc32/inc4_6/n1069 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_6/U10  ( .ZN(\ALUSHT/ALU/pkincout[27] ), 
        .A(\ALUSHT/ALU/pkincin[27] ), .B(\ALUSHT/ALU/inc32/inc4_6/n1071 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_6/U11  ( .Z(\ALUSHT/ALU/pkincout[26] ), 
        .A(\ALUSHT/ALU/pkincin[26] ), .B(\ALUSHT/ALU/inc32/inc4_6/n1070 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_7/U7  ( .Z(
        \ALUSHT/ALU/inc32/inc4_7/gp_out ), .A(\ALUSHT/ALU/pkincin[31] ), .B(
        \ALUSHT/ALU/pkincin[28] ), .C(\ALUSHT/ALU/pkincin[29] ), .D(
        \ALUSHT/ALU/pkincin[30] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_7/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_7/n1066 ), .A(\ALUSHT/ALU/pkincin[28] ), .B(
        \ALUSHT/ALU/inc32/gg_out[6] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_7/U13  ( .Z(\ALUSHT/ALU/pkincout[28] ), 
        .A(\ALUSHT/ALU/pkincin[28] ), .B(\ALUSHT/ALU/inc32/gg_out[6] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_7/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_7/n1068 ), .A(\ALUSHT/ALU/pkincin[30] ), .B(
        \ALUSHT/ALU/inc32/inc4_7/n1067 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_7/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_7/n1067 ), .A(\ALUSHT/ALU/inc32/inc4_7/n1066 ), 
        .B(\ALUSHT/ALU/pkincin[29] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_7/U12  ( .ZN(\ALUSHT/ALU/pkincout[29] ), 
        .A(\ALUSHT/ALU/pkincin[29] ), .B(\ALUSHT/ALU/inc32/inc4_7/n1066 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_7/U10  ( .ZN(\ALUSHT/ALU/pkincout[31] ), 
        .A(\ALUSHT/ALU/pkincin[31] ), .B(\ALUSHT/ALU/inc32/inc4_7/n1068 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_7/U11  ( .Z(\ALUSHT/ALU/pkincout[30] ), 
        .A(\ALUSHT/ALU/pkincin[30] ), .B(\ALUSHT/ALU/inc32/inc4_7/n1067 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_2/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[2] 
        ), .A(\ALUSHT/ALU/pkincin[11] ), .B(\ALUSHT/ALU/pkincin[8] ), .C(
        \ALUSHT/ALU/pkincin[9] ), .D(\ALUSHT/ALU/pkincin[10] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_2/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_2/n1063 ), .A(\ALUSHT/ALU/pkincin[8] ), .B(
        \ALUSHT/ALU/inc32/gg_out[1] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_2/U13  ( .Z(\ALUSHT/ALU/pkincout[8] ), 
        .A(\ALUSHT/ALU/pkincin[8] ), .B(\ALUSHT/ALU/inc32/gg_out[1] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_2/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_2/n1065 ), .A(\ALUSHT/ALU/pkincin[10] ), .B(
        \ALUSHT/ALU/inc32/inc4_2/n1064 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_2/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_2/n1064 ), .A(\ALUSHT/ALU/inc32/inc4_2/n1063 ), 
        .B(\ALUSHT/ALU/pkincin[9] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_2/U12  ( .ZN(\ALUSHT/ALU/pkincout[9] ), 
        .A(\ALUSHT/ALU/pkincin[9] ), .B(\ALUSHT/ALU/inc32/inc4_2/n1063 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_2/U10  ( .ZN(\ALUSHT/ALU/pkincout[11] ), 
        .A(\ALUSHT/ALU/pkincin[11] ), .B(\ALUSHT/ALU/inc32/inc4_2/n1065 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_2/U11  ( .Z(\ALUSHT/ALU/pkincout[10] ), 
        .A(\ALUSHT/ALU/pkincin[10] ), .B(\ALUSHT/ALU/inc32/inc4_2/n1064 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_3/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[3] 
        ), .A(\ALUSHT/ALU/pkincin[15] ), .B(\ALUSHT/ALU/pkincin[12] ), .C(
        \ALUSHT/ALU/pkincin[13] ), .D(\ALUSHT/ALU/pkincin[14] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_3/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_3/n1060 ), .A(\ALUSHT/ALU/pkincin[12] ), .B(
        \ALUSHT/ALU/inc32/gg_out[2] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_3/U13  ( .Z(\ALUSHT/ALU/pkincout[12] ), 
        .A(\ALUSHT/ALU/pkincin[12] ), .B(\ALUSHT/ALU/inc32/gg_out[2] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_3/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_3/n1062 ), .A(\ALUSHT/ALU/pkincin[14] ), .B(
        \ALUSHT/ALU/inc32/inc4_3/n1061 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_3/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_3/n1061 ), .A(\ALUSHT/ALU/inc32/inc4_3/n1060 ), 
        .B(\ALUSHT/ALU/pkincin[13] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_3/U12  ( .ZN(\ALUSHT/ALU/pkincout[13] ), 
        .A(\ALUSHT/ALU/pkincin[13] ), .B(\ALUSHT/ALU/inc32/inc4_3/n1060 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_3/U10  ( .ZN(\ALUSHT/ALU/pkincout[15] ), 
        .A(\ALUSHT/ALU/pkincin[15] ), .B(\ALUSHT/ALU/inc32/inc4_3/n1062 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_3/U11  ( .Z(\ALUSHT/ALU/pkincout[14] ), 
        .A(\ALUSHT/ALU/pkincin[14] ), .B(\ALUSHT/ALU/inc32/inc4_3/n1061 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_4/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[4] 
        ), .A(\ALUSHT/ALU/pkincin[19] ), .B(\ALUSHT/ALU/pkincin[16] ), .C(
        \ALUSHT/ALU/pkincin[17] ), .D(\ALUSHT/ALU/pkincin[18] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_4/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_4/n1057 ), .A(\ALUSHT/ALU/pkincin[16] ), .B(
        \ALUSHT/ALU/inc32/gg_out[3] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_4/U13  ( .Z(\ALUSHT/ALU/pkincout[16] ), 
        .A(\ALUSHT/ALU/pkincin[16] ), .B(\ALUSHT/ALU/inc32/gg_out[3] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_4/U14  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_4/n1059 ), .A(\ALUSHT/ALU/pkincin[18] ), .B(
        \ALUSHT/ALU/inc32/inc4_4/n1058 ) );
    snl_and12x1 \ALUSHT/ALU/inc32/inc4_4/U9  ( .Z(
        \ALUSHT/ALU/inc32/inc4_4/n1058 ), .A(\ALUSHT/ALU/inc32/inc4_4/n1057 ), 
        .B(\ALUSHT/ALU/pkincin[17] ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_4/U12  ( .ZN(\ALUSHT/ALU/pkincout[17] ), 
        .A(\ALUSHT/ALU/pkincin[17] ), .B(\ALUSHT/ALU/inc32/inc4_4/n1057 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_4/U10  ( .ZN(\ALUSHT/ALU/pkincout[19] ), 
        .A(\ALUSHT/ALU/pkincin[19] ), .B(\ALUSHT/ALU/inc32/inc4_4/n1059 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_4/U11  ( .Z(\ALUSHT/ALU/pkincout[18] ), 
        .A(\ALUSHT/ALU/pkincin[18] ), .B(\ALUSHT/ALU/inc32/inc4_4/n1058 ) );
    snl_and04x1 \ALUSHT/ALU/inc32/inc4_5/U7  ( .Z(\ALUSHT/ALU/inc32/gp_out[5] 
        ), .A(\ALUSHT/ALU/pkincin[23] ), .B(\ALUSHT/ALU/pkincin[20] ), .C(
        \ALUSHT/ALU/pkincin[21] ), .D(\ALUSHT/ALU/pkincin[22] ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_5/U8  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_5/n1052 ), .A(\ALUSHT/ALU/pkincin[20] ), .B(
        \ALUSHT/ALU/inc32/gg_out[4] ) );
    snl_aoi022x1 \ALUSHT/ALU/inc32/inc4_5/U13  ( .ZN(\ALUSHT/ALU/pkincout[21] 
        ), .A(\ALUSHT/ALU/pkincin[21] ), .B(\ALUSHT/ALU/inc32/inc4_5/n1056 ), 
        .C(\ALUSHT/ALU/inc32/inc4_5/n1053 ), .D(
        \ALUSHT/ALU/inc32/inc4_5/n1052 ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_5/U14  ( .Z(\ALUSHT/ALU/pkincout[20] ), 
        .A(\ALUSHT/ALU/pkincin[20] ), .B(\ALUSHT/ALU/inc32/gg_out[4] ) );
    snl_invx05 \ALUSHT/ALU/inc32/inc4_5/U9  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_5/n1053 ), .A(\ALUSHT/ALU/pkincin[21] ) );
    snl_xor2x0 \ALUSHT/ALU/inc32/inc4_5/U12  ( .Z(\ALUSHT/ALU/pkincout[22] ), 
        .A(\ALUSHT/ALU/pkincin[22] ), .B(\ALUSHT/ALU/inc32/inc4_5/n1054 ) );
    snl_nor02x1 \ALUSHT/ALU/inc32/inc4_5/U10  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_5/n1054 ), .A(\ALUSHT/ALU/inc32/inc4_5/n1053 ), 
        .B(\ALUSHT/ALU/inc32/inc4_5/n1052 ) );
    snl_nand02x1 \ALUSHT/ALU/inc32/inc4_5/U15  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_5/n1055 ), .A(\ALUSHT/ALU/pkincin[22] ), .B(
        \ALUSHT/ALU/inc32/inc4_5/n1054 ) );
    snl_xnor2x0 \ALUSHT/ALU/inc32/inc4_5/U11  ( .ZN(\ALUSHT/ALU/pkincout[23] ), 
        .A(\ALUSHT/ALU/pkincin[23] ), .B(\ALUSHT/ALU/inc32/inc4_5/n1055 ) );
    snl_invx05 \ALUSHT/ALU/inc32/inc4_5/U16  ( .ZN(
        \ALUSHT/ALU/inc32/inc4_5/n1056 ), .A(\ALUSHT/ALU/inc32/inc4_5/n1052 )
         );
endmodule

